// ----------------------------
// AXI to SRAM Adapter
// ----------------------------
// Author: Florian Zaruba (zarubaf@iis.ee.ethz.ch)
//
// Description: Manages AXI transactions
//              Supports all burst accesses but only on aligned addresses and with full data width.
//              Assertions should guide you if there is something unsupported happening.
//
module axi_mem_if #(
    parameter int unsigned AXI_ID_WIDTH      = 7,
    parameter int unsigned AXI_ADDR_WIDTH    = 48,
    parameter int unsigned AXI_DATA_WIDTH    = 128,
    parameter int unsigned AXI_USER_WIDTH    = 2
)(
    input    logic                        clk_i,    // Clock
    input    logic                        rst_ni,   // Asynchronous reset active low

    // AXI slave 
    input    logic                        aw_valid,
    output   logic                        aw_ready,
    input    logic [AXI_ADDR_WIDTH-1:0]   aw_addr,
    input    logic [AXI_ID_WIDTH-1  :0]   aw_id,
    input    logic [7:0]                  aw_len,
    input    logic [2:0]                  aw_size,
    input    logic [1:0]                  aw_burst,
    input    logic [3:0]                  aw_cache,
    input    logic [2:0]                  aw_prot,
    input    logic                        w_valid,
    output   logic                        w_ready,
    input    logic [AXI_DATA_WIDTH-1:0]   w_data,
    input    logic [15:0]                 w_strb,
    input    logic                        w_last,
    output   logic                        b_valid,
    input    logic                        b_ready,
    output   logic [AXI_ID_WIDTH-1  :0]   b_id,
    output   logic [1:0]                  b_resp,
    input    logic                        ar_valid,
    output   logic                        ar_ready,
    input    logic [AXI_ADDR_WIDTH-1:0]   ar_addr,
    input    logic [AXI_ID_WIDTH-1  :0]   ar_id,
    input    logic [7:0]                  ar_len,
    input    logic [2:0]                  ar_size,
    input    logic [1:0]                  ar_burst,
    input    logic [3:0]                  ar_cache,
    input    logic [2:0]                  ar_prot,
    output   logic                        r_valid,
    input    logic                        r_ready,
    output   logic [AXI_DATA_WIDTH-1:0]   r_data,
    output   logic [AXI_ID_WIDTH-1:0]     r_id,
    output   logic [1:0]                  r_resp,
    output   logic                        r_last,

    /// slave ram
    output   logic                        req_o,
    output   logic                        we_o,
    output   logic [AXI_ADDR_WIDTH-1:0]   addr_o,
    output   logic [AXI_DATA_WIDTH/8-1:0] be_o,
    output   logic [AXI_DATA_WIDTH-1:0]   data_o,
    input    logic [AXI_DATA_WIDTH-1:0]   data_i
);

    // AXI has the following rules governing the use of bursts:
    // - for wrapping bursts, the burst length must be 2, 4, 8, or 16
    // - a burst must not cross a 4KB address boundary
    // - early termination of bursts is not supported.
    typedef enum logic [1:0] { FIXED = 2'b00, INCR = 2'b01, WRAP = 2'b10} axi_burst_t;

    localparam LOG_NR_BYTES = $clog2(AXI_DATA_WIDTH/8);

    typedef struct packed {
        logic [AXI_ID_WIDTH-1:0]   id;
        logic [AXI_ADDR_WIDTH-1:0] addr;
        logic [7:0]                len;
        logic [2:0]                size;
        axi_burst_t                burst;
    } ax_req_t;

    // Registers
    enum logic [2:0] { IDLE, READ, WRITE, SEND_B, WAIT_WVALID }  state_d, state_q;
    ax_req_t                   ax_req_d, ax_req_q;
    logic [AXI_ADDR_WIDTH-1:0] req_addr_d, req_addr_q;
    logic [7:0]                cnt_d, cnt_q;

    function automatic logic [AXI_ADDR_WIDTH-1:0] get_wrap_boundary (input logic [AXI_ADDR_WIDTH-1:0] unaligned_address, input logic [7:0] len);
        logic [AXI_ADDR_WIDTH-1:0] warp_address = '0;
        //  for wrapping transfers ax_len can only be of size 1, 3, 7 or 15
        if (len == 4'b1)
            warp_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES];
        else if (len == 4'b11)
            warp_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES];
        else if (len == 4'b111)
            warp_address[AXI_ADDR_WIDTH-1:3+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:2+LOG_NR_BYTES];
        else if (len == 4'b1111)
            warp_address[AXI_ADDR_WIDTH-1:4+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:4+LOG_NR_BYTES];

        return warp_address;
    endfunction

    logic [AXI_ADDR_WIDTH-1:0] aligned_address;
    logic [AXI_ADDR_WIDTH-1:0] wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] upper_wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] cons_addr;

    always_comb begin
        // address generation
        aligned_address = {ax_req_q.addr[AXI_ADDR_WIDTH-1:LOG_NR_BYTES], {{LOG_NR_BYTES}{1'b0}}};
        wrap_boundary = get_wrap_boundary(ax_req_q.addr, ax_req_q.len);
        // this will overflow
        upper_wrap_boundary = wrap_boundary + ((ax_req_q.len + 1) << LOG_NR_BYTES);
        // calculate consecutive address
        cons_addr = aligned_address + (cnt_q << LOG_NR_BYTES);

        // Transaction attributes
        // default assignments
        state_d    = state_q;
        ax_req_d   = ax_req_q;
        req_addr_d = req_addr_q;
        cnt_d      = cnt_q;
        // Memory default assignments
        data_o = w_data;
        // user_o = w_user;
        be_o   = w_strb;
        we_o   = 1'b0;
        req_o  = 1'b0;
        addr_o = '0;
        // AXI assignments
        // request
        aw_ready = 1'b0;
        ar_ready = 1'b0;
        // read response channel
        r_valid  = 1'b0;
        r_data   = data_i;
        r_resp   = '0;
        r_last   = '0;
        r_id     = ax_req_q.id;
        // r_user   = user_i;
        // slave write data channel
        w_ready  = 1'b0;
        // write response channel
        b_valid  = 1'b0;
        b_resp   = 1'b0;
        b_id     = 1'b0;
        // b_user   = 1'b0;

        case (state_q)

            IDLE: begin
                // Wait for a read or write
                // ------------
                // Read
                // ------------
                if (ar_valid) begin
                    ar_ready = 1'b1;
                    // sample ax
                    ax_req_d       = {ar_id, ar_addr, ar_len, ar_size, ar_burst};
                    state_d        = READ;
                    //  we can request the first address, this saves us time
                    req_o          = 1'b1;
                    addr_o         = ar_addr;
                    // save the address
                    req_addr_d     = ar_addr;
                    // save the ar_len
                    cnt_d          = 1;
                // ------------
                // Write
                // ------------
                end else if (aw_valid) begin
                    aw_ready = 1'b1;
                    w_ready  = 1'b1;
                    addr_o         = aw_addr;
                    // sample ax
                    ax_req_d       = {aw_id, aw_addr, aw_len, aw_size, aw_burst};
                    // we've got our first w_valid so start the write process
                    if (w_valid) begin
                        req_o          = 1'b1;
                        we_o           = 1'b1;
                        state_d        = (w_last) ? SEND_B : WRITE;
                        cnt_d          = 1;
                    // we still have to wait for the first w_valid to arrive
                    end else
                        state_d = WAIT_WVALID;
                end
            end

            // ~> we are still missing a w_valid
            WAIT_WVALID: begin
                w_ready = 1'b1;
                addr_o = ax_req_q.addr;
                // we can now make our first request
                if (w_valid) begin
                    req_o          = 1'b1;
                    we_o           = 1'b1;
                    state_d        = (w_last) ? SEND_B : WRITE;
                    cnt_d          = 1;
                end
            end

            READ: begin
                // keep request to memory high
                req_o  = 1'b1;
                addr_o = req_addr_q;
                // send the response
                r_valid = 1'b1;
                r_data  = data_i;
                // r_user  = user_i;
                r_id    = ax_req_q.id;
                r_last  = (cnt_q == ax_req_q.len + 1);

                // check that the master is ready, the slave must not wait on this
                if (r_ready) begin
                    // ----------------------------
                    // Next address generation
                    // ----------------------------
                    // handle the correct burst type
                    case (ax_req_q.burst)
                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            // check if the address reached warp boundary
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            // address warped beyond boundary
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len - 1) << LOG_NR_BYTES);
                            // we are still in the incremental regime
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    // we need to change the address here for the upcoming request
                    // we sent the last byte -> go back to idle
                    if (r_last) begin
                        state_d = IDLE;
                        // we already got everything
                        req_o = 1'b0;
                    end
                    // save the request address for the next cycle
                    req_addr_d = addr_o;
                    // we can decrease the counter as the master has consumed the read data
                    cnt_d = cnt_q + 1;
                    // TODO: configure correct byte-lane
                end
            end
            // ~> we already wrote the first word here
            WRITE: begin

                w_ready = 1'b1;

                // consume a word here
                if (w_valid) begin
                    req_o         = 1'b1;
                    we_o          = 1'b1;
                    // ----------------------------
                    // Next address generation
                    // ----------------------------
                    // handle the correct burst type
                    case (ax_req_q.burst)

                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            // check if the address reached warp boundary
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            // address warped beyond boundary
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len - 1) << LOG_NR_BYTES);
                            // we are still in the incremental regime
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    // save the request address for the next cycle
                    req_addr_d = addr_o;
                    // we can decrease the counter as the master has consumed the read data
                    cnt_d = cnt_q + 1;

                    if (w_last)
                        state_d = SEND_B;
                end
            end
            // ~> send a write acknowledge back
            SEND_B: begin
                b_valid = 1'b1;
                b_id    = ax_req_q.id;
                if (b_ready)
                    state_d = IDLE;
            end

        endcase
    end
    // --------------
    // Registers
    // --------------
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q    <= IDLE;
            ax_req_q  <= '0;
            req_addr_q <= '0;
            cnt_q      <= '0;
        end else begin
            state_q    <= state_d;
            ax_req_q   <= ax_req_d;
            req_addr_q <= req_addr_d;
            cnt_q      <= cnt_d;
        end
    end
endmodule


