/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @23
module aq_vfmau_lza_double (
  // &Ports, @24
  input    wire  [110:0]  addend,
  input    wire           sub_vld,
  input    wire  [110:0]  summand,
  input    wire  [110:0]  upper_limit,
  output   reg   [6  :0]  lza_result
); 



// &Regs; @25

// &Wires; @26
wire    [110:0]  carry_d;     
wire    [110:0]  carry_g;     
wire    [110:0]  carry_p;     
wire    [110:0]  data_for_ff1; 
wire    [110:0]  lza_precod;  


parameter DATA_WIDTH   = 111;
parameter DATA_WIDTH_D = 111;
parameter DATA_WIDTH_S = 53;

// &CombBeg; @81
// &CombEnd; @144
// &CombBeg; @174
// &CombEnd; @232
 //==========================================================
//                   Signal Pre-encode
//==========================================================
//----------------------------------------------------------
//                   Signal preparation
//----------------------------------------------------------
// carry_p: carry propagete
// carry_g: carry generate
// carry_d: carry delete
assign carry_p[DATA_WIDTH-1:0] =   summand[DATA_WIDTH-1:0] ^ addend[DATA_WIDTH-1:0];
assign carry_g[DATA_WIDTH-1:0] =   summand[DATA_WIDTH-1:0] & addend[DATA_WIDTH-1:0];
assign carry_d[DATA_WIDTH-1:0] = ~(summand[DATA_WIDTH-1:0] | addend[DATA_WIDTH-1:0]);
//----------------------------------------------------------
//                   Signal decode
//----------------------------------------------------------
//pre-predecode for leading zero anticipation
assign lza_precod[0] = 
     carry_p[1] && (carry_g[0] && sub_vld || carry_d[0])
 || !carry_p[1] && (carry_d[0] && sub_vld || carry_g[0]);

assign lza_precod[DATA_WIDTH-1] = 
     sub_vld && (carry_g[DATA_WIDTH-1] && !carry_d[DATA_WIDTH-2] 
 ||  carry_d[DATA_WIDTH-1] && !carry_g[DATA_WIDTH-2])
 || !sub_vld && (carry_d[DATA_WIDTH-1] && !carry_d[DATA_WIDTH-2] 
 || !carry_d[DATA_WIDTH-1]);

assign lza_precod[DATA_WIDTH-2:1] = 
    carry_p[DATA_WIDTH-1:2] & (carry_g[DATA_WIDTH-2:1] & ~carry_d[DATA_WIDTH-3:0] 
 |  carry_d[DATA_WIDTH-2:1] & ~carry_g[DATA_WIDTH-3:0])
 | ~carry_p[DATA_WIDTH-1:2] & (carry_g[DATA_WIDTH-2:1] & ~carry_g[DATA_WIDTH-3:0] 
 |  carry_d[DATA_WIDTH-2:1] & ~carry_d[DATA_WIDTH-3:0]);


//==========================================================
//                     LZA coding
//==========================================================
assign data_for_ff1[DATA_WIDTH-1:0] = lza_precod[DATA_WIDTH-1:0] | upper_limit[DATA_WIDTH-1:0];
// &CombBeg; @276
always @( data_for_ff1[110:0])
begin
casez(data_for_ff1[DATA_WIDTH-1:0])
  111'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd0;
  111'b01?????????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd1;
  111'b001????????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd2;
  111'b0001???????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd3;
  111'b00001??????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd4;
  111'b000001?????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd5;
  111'b0000001????????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd6;
  111'b00000001???????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd7;
  111'b000000001??????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd8;
  111'b0000000001?????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd9;
  111'b00000000001????????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd10;
  111'b000000000001???????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd11;
  111'b0000000000001??????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd12;
  111'b00000000000001?????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd13;
  111'b000000000000001????????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd14;
  111'b0000000000000001???????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd15;
  111'b00000000000000001??????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd16;
  111'b000000000000000001?????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd17;
  111'b0000000000000000001????????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd18;
  111'b00000000000000000001???????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd19;
  111'b000000000000000000001??????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd20;
  111'b0000000000000000000001?????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd21;
  111'b00000000000000000000001????????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd22;
  111'b000000000000000000000001???????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd23;
  111'b0000000000000000000000001??????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd24;
  111'b00000000000000000000000001?????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd25;
  111'b000000000000000000000000001????????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd26;
  111'b0000000000000000000000000001???????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd27;
  111'b00000000000000000000000000001??????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd28;
  111'b000000000000000000000000000001?????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd29;
  111'b0000000000000000000000000000001????????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd30;
  111'b00000000000000000000000000000001???????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd31;
  111'b000000000000000000000000000000001??????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd32;
  111'b0000000000000000000000000000000001?????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd33;
  111'b00000000000000000000000000000000001????????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd34;
  111'b000000000000000000000000000000000001???????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd35;
  111'b0000000000000000000000000000000000001??????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd36;
  111'b00000000000000000000000000000000000001?????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd37;
  111'b000000000000000000000000000000000000001????????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd38;
  111'b0000000000000000000000000000000000000001???????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd39;
  111'b00000000000000000000000000000000000000001??????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd40;
  111'b000000000000000000000000000000000000000001?????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd41;
  111'b0000000000000000000000000000000000000000001????????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd42;
  111'b00000000000000000000000000000000000000000001???????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd43;
  111'b000000000000000000000000000000000000000000001??????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd44;
  111'b0000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd45;
  111'b00000000000000000000000000000000000000000000001????????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd46;
  111'b000000000000000000000000000000000000000000000001???????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd47;
  111'b0000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd48;
  111'b00000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd49;
  111'b000000000000000000000000000000000000000000000000001????????????????????????????????????????????????????????????:lza_result[6:0] = 7'd50;
  111'b0000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????????????:lza_result[6:0] = 7'd51;
  111'b00000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????????:lza_result[6:0] = 7'd52;
  111'b000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????:lza_result[6:0] = 7'd53;
  111'b0000000000000000000000000000000000000000000000000000001????????????????????????????????????????????????????????:lza_result[6:0] = 7'd54;
  111'b00000000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????????:lza_result[6:0] = 7'd55;
  111'b000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????:lza_result[6:0] = 7'd56;
  111'b0000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????:lza_result[6:0] = 7'd57;
  111'b00000000000000000000000000000000000000000000000000000000001????????????????????????????????????????????????????:lza_result[6:0] = 7'd58;
  111'b000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????:lza_result[6:0] = 7'd59;
  111'b0000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????:lza_result[6:0] = 7'd60;
  111'b00000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????:lza_result[6:0] = 7'd61;
  111'b000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????????????????:lza_result[6:0] = 7'd62;
  111'b0000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????????????:lza_result[6:0] = 7'd63;
  111'b00000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????????:lza_result[6:0] = 7'd64;
  111'b000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????:lza_result[6:0] = 7'd65;
  111'b0000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????????????:lza_result[6:0] = 7'd66;
  111'b00000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????????:lza_result[6:0] = 7'd67;
  111'b000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????:lza_result[6:0] = 7'd68;
  111'b0000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????:lza_result[6:0] = 7'd69;
  111'b00000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????????:lza_result[6:0] = 7'd70;
  111'b000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????:lza_result[6:0] = 7'd71;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????:lza_result[6:0] = 7'd72;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????:lza_result[6:0] = 7'd73;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????:lza_result[6:0] = 7'd74;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????:lza_result[6:0] = 7'd75;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????:lza_result[6:0] = 7'd76;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????:lza_result[6:0] = 7'd77;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????:lza_result[6:0] = 7'd78;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????:lza_result[6:0] = 7'd79;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????:lza_result[6:0] = 7'd80;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????:lza_result[6:0] = 7'd81;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????:lza_result[6:0] = 7'd82;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????:lza_result[6:0] = 7'd83;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????:lza_result[6:0] = 7'd84;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????:lza_result[6:0] = 7'd85;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????:lza_result[6:0] = 7'd86;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????:lza_result[6:0] = 7'd87;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????:lza_result[6:0] = 7'd88;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????:lza_result[6:0] = 7'd89;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????:lza_result[6:0] = 7'd90;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????:lza_result[6:0] = 7'd91;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????:lza_result[6:0] = 7'd92;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????:lza_result[6:0] = 7'd93;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????:lza_result[6:0] = 7'd94;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????:lza_result[6:0] = 7'd95;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????:lza_result[6:0] = 7'd96;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????:lza_result[6:0] = 7'd97;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????:lza_result[6:0] = 7'd98;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????:lza_result[6:0] = 7'd99;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????:lza_result[6:0] = 7'd100;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????:lza_result[6:0] = 7'd101;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????:lza_result[6:0] = 7'd102;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????:lza_result[6:0] = 7'd103;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????:lza_result[6:0] = 7'd104;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????:lza_result[6:0] = 7'd105;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????:lza_result[6:0] = 7'd106;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???:lza_result[6:0] = 7'd107;
  111'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??:lza_result[6:0] = 7'd108;
  111'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?:lza_result[6:0] = 7'd109;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001:lza_result[6:0] = 7'd110;
  111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:lza_result[6:0] = 7'd111;
  default                                                                                                             :lza_result[6:0] = 7'd0;
endcase
// &CombEnd; @392
end


// &ModuleEnd; @396
endmodule



