/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/
module ct_cp0_top (
  // &Ports, @25
  input    wire  [39 :0]  biu_cp0_apb_base,
  input    wire           biu_cp0_cmplt,
  input    wire  [2  :0]  biu_cp0_coreid,
  input    wire  [7  :0]  ext_interrupt,
  input    wire           biu_cp0_me_int,
  input    wire           biu_cp0_ms_int,
  input    wire           biu_cp0_mt_int,
  input    wire  [127:0]  biu_cp0_rdata,
  input    wire  [39 :0]  biu_cp0_rvba,
  input    wire           biu_cp0_se_int,
  input    wire           biu_cp0_ss_int,
  input    wire           biu_cp0_st_int,
  input    wire           biu_yy_xx_no_op,
  input    wire           cpurst_b,
  input    wire           forever_cpuclk,
  input    wire           had_cp0_xx_dbg,
  input    wire           hpcp_cp0_cmplt,
  input    wire  [63 :0]  hpcp_cp0_data,
  input    wire           hpcp_cp0_int_vld,
  input    wire           hpcp_cp0_sce,
  input    wire  [6  :0]  idu_cp0_fesr_acc_updt_val,
  input    wire           idu_cp0_fesr_acc_updt_vld,
  input    wire  [4  :0]  idu_cp0_rf_func,
  input    wire           idu_cp0_rf_gateclk_sel,
  input    wire  [6  :0]  idu_cp0_rf_iid,
  input    wire  [31 :0]  idu_cp0_rf_opcode,
  input    wire  [6  :0]  idu_cp0_rf_preg,
  input    wire           idu_cp0_rf_sel,
  input    wire  [63 :0]  idu_cp0_rf_src0,
  input    wire  [63 :0]  idu_cp0_rf_src1,
  input    wire           ifu_cp0_bht_inv_done,
  input    wire           ifu_cp0_btb_inv_done,
  input    wire           ifu_cp0_icache_inv_done,
  input    wire  [127:0]  ifu_cp0_icache_read_data,
  input    wire           ifu_cp0_icache_read_data_vld,
  input    wire           ifu_cp0_ind_btb_inv_done,
  input    wire           ifu_cp0_rst_inv_req,
  input    wire           ifu_yy_xx_no_op,
  input    wire           lsu_cp0_dcache_done,
  input    wire  [127:0]  lsu_cp0_dcache_read_data,
  input    wire           lsu_cp0_dcache_read_data_vld,
  input    wire  [63 :0]  lsu_cp0_ld_va,
  input    wire  [39 :0]  lsu_cp0_ld_pa,
  input    wire           lsu_cp0_ld_vld,
  input    wire           lsu_yy_xx_no_op,
  input    wire           mmu_cp0_cmplt,
  input    wire  [63 :0]  mmu_cp0_data,
  input    wire  [63 :0]  mmu_cp0_satp_data,
  input    wire           mmu_cp0_tlb_done,
  input    wire           mmu_cp0_type,
  input    wire  [26 :0]  mmu_cp0_vpn,
  input    wire           mmu_cp0_fst_vld,
  input    wire  [39 :0]  mmu_cp0_fst_addr,
  input    wire           mmu_cp0_scd_vld,
  input    wire  [39 :0]  mmu_cp0_scd_addr,
  input    wire           mmu_cp0_thd_vld,
  input    wire  [39 :0]  mmu_cp0_thd_addr,
  input    wire           mmu_yy_xx_no_op,
  input    wire           pad_yy_icg_scan_en,
  input    wire  [63 :0]  pmp_cp0_data,
  input    wire  [63 :0]  rtu_cp0_epc,
  input    wire           rtu_cp0_expt_gateclk_vld,
  input    wire  [63 :0]  rtu_cp0_expt_mtval,
  input    wire           rtu_cp0_expt_vld,
  input    wire           rtu_cp0_fp_dirty_vld,
  input    wire           rtu_cp0_int_ack,
  input    wire           rtu_cp0_vec_dirty_vld,
  input    wire           rtu_cp0_vsetvl_vill,
  input    wire  [7  :0]  rtu_cp0_vsetvl_vl,
  input    wire           rtu_cp0_vsetvl_vl_vld,
  input    wire  [1  :0]  rtu_cp0_vsetvl_vlmul,
  input    wire  [2  :0]  rtu_cp0_vsetvl_vsew,
  input    wire           rtu_cp0_vsetvl_vtype_vld,
  input    wire  [6  :0]  rtu_cp0_vstart,
  input    wire           rtu_cp0_vstart_vld,
  input    wire           rtu_yy_xx_commit0,
  input    wire  [6  :0]  rtu_yy_xx_commit0_iid,
  input    wire           rtu_yy_xx_dbgon,
  input    wire  [15 :0]  rtu_yy_xx_expt_vec,
  input    wire           rtu_yy_xx_flush,
  input    wire  [63 :0]  sysio_core_gl_stable_timer,
  input    wire           sysio_core_restart_vld,
  input    wire           core_sysio_restart_grnt,
  input    wire           sysio_core_cp0_update_ipi_status_en,
  input    wire  [31 :0]  sysio_core_cp0_update_ipi_status_src,
  input    wire           sysio_core_cp0_update_mailbox0_en,
  input    wire           sysio_core_cp0_update_mailbox1_en,
  input    wire           sysio_core_cp0_update_mailbox2_en,
  input    wire           sysio_core_cp0_update_mailbox3_en,
  input    wire           sysio_core_cp0_req_grnt,
  input    wire  [3  :0]  sysio_core_cp0_update_bit_sel,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_src0,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_src1,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_src2,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_src3,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_mask0,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_mask1,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_mask2,
  input    wire  [31 :0]  sysio_core_cp0_update_mailbox_mask3,
  output   wire           cp0_biu_icg_en,
  output   wire  [1  :0]  cp0_biu_lpmd_b,
  output   wire  [15 :0]  cp0_biu_op,
  output   wire           cp0_biu_sel,
  output   wire  [63 :0]  cp0_biu_wdata,
  output   wire  [31 :0]  cp0_had_cpuid_0,
  output   wire  [3  :0]  cp0_had_debug_info,
  output   wire  [1  :0]  cp0_had_lpmd_b,
  output   wire  [1  :0]  cp0_had_trace_pm_wdata,
  output   wire           cp0_had_trace_pm_wen,
  output   wire           cp0_hpcp_icg_en,
  output   wire  [11 :0]  cp0_hpcp_index,
  output   wire           cp0_hpcp_int_disable,
  output   wire  [31 :0]  cp0_hpcp_mcntwen,
  output   wire  [3  :0]  cp0_hpcp_op,
  output   wire           cp0_hpcp_pmdm,
  output   wire           cp0_hpcp_pmds,
  output   wire           cp0_hpcp_pmdu,
  output   wire           cp0_hpcp_sel,
  output   wire  [63 :0]  cp0_hpcp_src0,
  output   wire  [63 :0]  cp0_hpcp_wdata,
  output   wire           cp0_idu_cskyee,
  output   wire           cp0_idu_dlb_disable,
  output   wire  [2  :0]  cp0_idu_frm,
  output   wire  [1  :0]  cp0_idu_fs,
  output   wire           cp0_idu_icg_en,
  output   wire           cp0_idu_iq_bypass_disable,
  output   wire           cp0_idu_rob_fold_disable,
  output   wire           cp0_idu_src2_fwd_disable,
  output   wire           cp0_idu_srcv2_fwd_disable,
  output   wire           cp0_idu_vill,
  output   wire  [1  :0]  cp0_idu_vs,
  output   wire  [6  :0]  cp0_idu_vstart,
  output   wire           cp0_idu_zero_delay_move_disable,
  output   wire           cp0_ifu_bht_en,
  output   wire           cp0_ifu_bht_inv,
  output   wire           cp0_ifu_btb_en,
  output   wire           cp0_ifu_btb_inv,
  output   wire           cp0_ifu_icache_en,
  output   wire           cp0_ifu_icache_inv,
  output   wire           cp0_ifu_icache_pref_en,
  output   wire  [16 :0]  cp0_ifu_icache_read_index,
  output   wire           cp0_ifu_icache_read_req,
  output   wire           cp0_ifu_icache_read_tag,
  output   wire           cp0_ifu_icache_read_way,
  output   wire           cp0_ifu_icg_en,
  output   wire           cp0_ifu_ind_btb_en,
  output   wire           cp0_ifu_ind_btb_inv,
  output   wire           cp0_ifu_insde,
  output   wire           cp0_ifu_iwpe,
  output   wire           cp0_ifu_l0btb_en,
  output   wire           cp0_ifu_lbuf_en,
  output   wire           cp0_ifu_no_op_req,
  output   wire           cp0_ifu_nsfe,
  output   wire           cp0_ifu_ras_en,
  output   wire           cp0_ifu_rst_inv_done,
  output   wire           cp0_ifu_boot_stall,
  output   wire  [39 :0]  cp0_ifu_rvbr,
  output   wire  [39 :0]  cp0_ifu_vbr,
  output   wire  [2  :0]  cp0_ifu_ecfg_vs,
  output   wire  [63 :0]  cp0_ifu_eentry,
  output   wire  [7  :0]  cp0_ifu_vl,
  output   wire  [1  :0]  cp0_ifu_vlmul,
  output   wire           cp0_ifu_vsetvli_pred_disable,
  output   wire           cp0_ifu_vsetvli_pred_mode,
  output   wire  [2  :0]  cp0_ifu_vsew,
  output   wire           cp0_iu_div_entry_disable,
  output   wire           cp0_iu_div_entry_disable_clr,
  output   wire           cp0_iu_ex3_abnormal,
  output   wire  [62 :0]  cp0_iu_ex3_efpc,
  output   wire           cp0_iu_ex3_efpc_vld,
  output   wire  [4  :0]  cp0_iu_ex3_expt_vec,
  output   wire           cp0_iu_ex3_expt_vld,
  output   wire           cp0_iu_ex3_flush,
  output   wire  [6  :0]  cp0_iu_ex3_iid,
  output   wire           cp0_iu_ex3_inst_vld,
  output   wire  [31 :0]  cp0_iu_ex3_mtval,
  output   wire  [63 :0]  cp0_iu_ex3_rslt_data,
  output   wire  [6  :0]  cp0_iu_ex3_rslt_preg,
  output   wire  [4  :0]  cp0_iu_ex3_rslt_dreg,
  output   wire           cp0_iu_ex3_rslt_vld,
  output   wire           cp0_iu_icg_en,
  output   wire           cp0_iu_bju_chflw_en,
  output   wire           cp0_iu_vill,
  output   wire  [7  :0]  cp0_iu_vl,
  output   wire           cp0_iu_vsetvli_pre_decd_disable,
  output   wire  [6  :0]  cp0_iu_vstart,
  output   wire  [63 :0]  cp0_iu_timer,
  output   wire           cp0_lsu_amr,
  output   wire           cp0_lsu_amr2,
  output   wire           cp0_lsu_cb_aclr_dis,
  output   wire           cp0_lsu_corr_dis,
  output   wire           cp0_lsu_ctc_flush_dis,
  output   wire           cp0_lsu_da_fwd_dis,
  output   wire           cp0_lsu_dcache_clr,
  output   wire           cp0_lsu_dcache_en,
  output   wire           cp0_lsu_dcache_inv,
  output   wire  [1  :0]  cp0_lsu_dcache_pref_dist,
  output   wire           cp0_lsu_dcache_pref_en,
  output   wire  [16 :0]  cp0_lsu_dcache_read_index,
  output   wire           cp0_lsu_dcache_read_ld_tag,
  output   wire           cp0_lsu_dcache_read_req,
  output   wire           cp0_lsu_dcache_read_st_tag,
  output   wire           cp0_lsu_dcache_read_way,
  output   wire           cp0_lsu_fencei_broad_dis,
  output   wire           cp0_lsu_fencerw_broad_dis,
  output   wire           cp0_lsu_icg_en,
  output   wire  [1  :0]  cp0_lsu_l2_pref_dist,
  output   wire           cp0_lsu_l2_pref_en,
  output   wire           cp0_lsu_l2_st_pref_en,
  output   wire           cp0_lsu_mm,
  output   wire           cp0_lsu_no_op_req,
  output   wire           cp0_lsu_nsfe,
  output   wire           cp0_lsu_pfu_mmu_dis,
  output   wire  [29 :0]  cp0_lsu_timeout_cnt,
  output   wire           cp0_lsu_tlb_broad_dis,
  output   wire           cp0_lsu_tvm,
  output   wire           cp0_lsu_ucme,
  output   wire  [6  :0]  cp0_lsu_vstart,
  output   wire           cp0_lsu_wa,
  output   wire           cp0_lsu_wr_burst_dis,
  output   wire           cp0_mmu_cskyee,
  output   wire           cp0_mmu_icg_en,
  output   wire           cp0_mmu_maee,
  output   wire  [1  :0]  cp0_mmu_mpp,
  output   wire           cp0_mmu_mprv,
  output   wire           cp0_mmu_mxr,
  output   wire           cp0_mmu_no_op_req,
  output   wire           cp0_mmu_ptw_en,
  output   wire  [1  :0]  cp0_mmu_reg_num,
  output   wire           cp0_mmu_satp_sel,
  output   wire           cp0_mmu_sum,
  output   wire           cp0_mmu_tlb_all_inv,
  output   wire  [63 :0]  cp0_mmu_wdata,
  output   wire           cp0_mmu_wreg,
  output   wire           cp0_mmu_crmd_da,
  output   wire           cp0_mmu_crmd_pg,
  output   wire  [15: 0]  cp0_mmu_cur_asid,
  output   wire  [1 : 0]  cp0_mmu_da_mode_datf,
  output   wire  [1 : 0]  cp0_mmu_da_mode_datm,
  output   wire  [63: 0]  cp0_mmu_ptw_pgdl,
  output   wire  [63: 0]  cp0_mmu_ptw_pgdh,
  output   wire  [63: 0]  cp0_mmu_dmw0,
  output   wire  [63: 0]  cp0_mmu_dmw1,
  output   wire  [63: 0]  cp0_mmu_dmw2,
  output   wire  [63: 0]  cp0_mmu_dmw3,
  output   wire  [63 :0]  cp0_pad_mstatus,
  output   wire           cp0_pmp_icg_en,
  output   wire  [1  :0]  cp0_pmp_mpp,
  output   wire           cp0_pmp_mprv,
  output   wire  [4  :0]  cp0_pmp_reg_num,
  output   wire  [63 :0]  cp0_pmp_wdata,
  output   wire           cp0_pmp_wreg,
  output   wire           cp0_rtu_icg_en,
  output   wire           cp0_rtu_srt_en,
  output   wire           cp0_rtu_xx_int_b,
  output   wire  [12 :0]  cp0_rtu_xx_vec,
  output   wire  [63 :0]  cp0_vfpu_fcsr,
  output   wire  [31 :0]  cp0_vfpu_fxcr,
  output   wire           cp0_vfpu_icg_en,
  output   wire  [7  :0]  cp0_vfpu_vl,
  output   wire           cp0_xx_core_arch,
  output   wire           cp0_xx_core_icg_en,
  output   wire           core_sysio_wr_req,
  output   wire  [3  :0]  core_sysio_wr_sel,
  output   wire  [31 :0]  core_sysio_wr_ipi_send_data,
  output   wire  [63 :0]  core_sysio_wr_mail_box_send_data,
  output   wire  [63 :0]  core_sysio_mailbox0_data,
  output   wire           cp0_yy_clk_en,
  output   wire           cp0_yy_dcache_pref_en,
  output   wire           cp0_yy_hyper,
  output   wire  [1  :0]  cp0_yy_priv_mode,
  output   wire           cp0_yy_virtual_mode
); 



// &Regs; @26
// &Wires; @27
wire             cp0_mret;                       
wire             cp0_ertn;                       
wire             cp0_cprs;                       
wire             cp0_sret;                       
wire             inst_lpmd_ex1_ex2;              
wire    [11 :0]  iui_regs_addr;                  
wire             iui_regs_csr_wr;                
wire             iui_regs_csrw;                  
wire             iui_regs_ex3_inst_csr;          
wire             iui_regs_inst_mret;             
wire             iui_regs_inst_ertn;             
wire             iui_regs_inst_sret;             
wire             iui_regs_inv_expt;              
wire    [31 :0]  iui_regs_opcode;                
wire    [63 :0]  iui_regs_ori_src0;              
wire    [63 :0]  iui_regs_cpu_cfg_code;              
wire             iui_regs_rst_inv_d;             
wire             iui_regs_rst_inv_i;             
wire             iui_regs_sel;                   
wire             iui_regs_sel_ipi;                   
wire    [63 :0]  iui_regs_src0;                  
wire    [1  :0]  iui_top_cur_state;              
wire             lpmd_cmplt;                     
wire    [1  :0]  lpmd_top_cur_state;             
wire             regs_iui_cfr_no_op;             
wire             regs_iui_chk_vld;               
wire             regs_iui_cindex_l2;             
wire             regs_iui_cins_no_op;            
wire             regs_iui_cskyee;                
wire    [63 :0]  regs_iui_data_out;              
wire    [63 :0]  regs_iui_iocsr_data_out;              
wire    [63 :0]  regs_iui_mailbox0_data;              
wire    [63 :0]  regs_iui_cfg_data_out;              
wire             regs_iui_dca_sel;               
wire             regs_iui_fs_off;                
wire             regs_iui_hpcp_regs_sel;         
wire             regs_iui_hpcp_scr_inv;          
wire    [14 :0]  regs_iui_int_sel;               
wire             regs_iui_l2_regs_sel;           
wire    [1  :0]  regs_iui_pm;                    
wire    [3  :0]  regs_iui_reg_idx;               
wire             regs_iui_scnt_inv;              
wire             regs_iui_tee_ff;                
wire             regs_iui_tee_vld;               
wire             regs_iui_tsr;                   
wire             regs_iui_tvm;                   
wire             regs_iui_tw;                    
wire             regs_iui_ucnt_inv;              
wire             regs_iui_v;                     
wire             regs_iui_vs_off;                
wire    [2  :0]  regs_iui_ecfg_vs;                
wire    [63 :0]  regs_iui_wdata;                 
wire             regs_lpmd_int_vld;              
wire             regs_xx_icg_en;                 
wire    [15 :0]  iui_regs_iocsr_addr;
wire    [63 :0]  iui_ipi_regs_src;
wire             iui_update_ipi_status_en;
wire    [31 :0]  iui_update_ipi_status_src;
wire             iui_update_ipi_mailbox0_en;
wire             iui_update_ipi_mailbox1_en;
wire             iui_update_ipi_mailbox2_en;
wire             iui_update_ipi_mailbox3_en;
wire    [ 3 :0]  iui_update_ipi_mailbox_sel;
wire    [31 :0]  iui_update_ipi_regs_src0;
wire    [31 :0]  iui_update_ipi_regs_src1;
wire    [31 :0]  iui_update_ipi_regs_src2;
wire    [31 :0]  iui_update_ipi_regs_src3;
wire    [31 :0]  iui_update_ipi_regs_mask0;
wire    [31 :0]  iui_update_ipi_regs_mask1;
wire    [31 :0]  iui_update_ipi_regs_mask2;
wire    [31 :0]  iui_update_ipi_regs_mask3;


// &Force ("output","cp0_yy_clk_en"); @30

// &Instance("ct_cp0_iui", "x_ct_cp0_iui"); @32
ct_cp0_iui x_ct_cp0_iui (
  .biu_cp0_cmplt                        (biu_cp0_cmplt                        ),
  .biu_cp0_rdata                        (biu_cp0_rdata                        ),
  .biu_cp0_coreid                       (biu_cp0_coreid                       ),
  .cp0_biu_op                           (cp0_biu_op                           ),
  .cp0_biu_sel                          (cp0_biu_sel                          ),
  .cp0_biu_wdata                        (cp0_biu_wdata                        ),
  .cp0_hpcp_op                          (cp0_hpcp_op                          ),
  .cp0_hpcp_sel                         (cp0_hpcp_sel                         ),
  .cp0_hpcp_src0                        (cp0_hpcp_src0                        ),
  .cp0_ifu_rst_inv_done                 (cp0_ifu_rst_inv_done                 ),
  .cp0_ifu_boot_stall                   (cp0_ifu_boot_stall                   ),
  .cp0_iu_ex3_abnormal                  (cp0_iu_ex3_abnormal                  ),
  .cp0_iu_ex3_expt_vec                  (cp0_iu_ex3_expt_vec                  ),
  .cp0_iu_ex3_expt_vld                  (cp0_iu_ex3_expt_vld                  ),
  .cp0_iu_ex3_flush                     (cp0_iu_ex3_flush                     ),
  .cp0_iu_ex3_iid                       (cp0_iu_ex3_iid                       ),
  .cp0_iu_ex3_inst_vld                  (cp0_iu_ex3_inst_vld                  ),
  .cp0_iu_ex3_mtval                     (cp0_iu_ex3_mtval                     ),
  .cp0_iu_ex3_rslt_data                 (cp0_iu_ex3_rslt_data                 ),
  .cp0_iu_ex3_rslt_preg                 (cp0_iu_ex3_rslt_preg                 ),
  .cp0_iu_ex3_rslt_dreg                 (cp0_iu_ex3_rslt_dreg                 ),
  .cp0_iu_ex3_rslt_vld                  (cp0_iu_ex3_rslt_vld                  ),
  .cp0_mmu_tlb_all_inv                  (cp0_mmu_tlb_all_inv                  ),
  .cp0_mret                             (cp0_mret                             ),
  .cp0_ertn                             (cp0_ertn                             ),
  .cp0_cprs                             (cp0_cprs                             ),
  .cp0_rtu_xx_int_b                     (cp0_rtu_xx_int_b                     ),
  .cp0_rtu_xx_vec                       (cp0_rtu_xx_vec                       ),
  .cp0_sret                             (cp0_sret                             ),
  .cp0_yy_clk_en                        (cp0_yy_clk_en                        ),
  .core_sysio_wr_req                    (core_sysio_wr_req                    ),
  .core_sysio_wr_sel                    (core_sysio_wr_sel                    ),
  .core_sysio_wr_ipi_send_data          (core_sysio_wr_ipi_send_data          ),
  .core_sysio_wr_mail_box_send_data     (core_sysio_wr_mail_box_send_data     ),
  .core_sysio_mailbox0_data             (core_sysio_mailbox0_data             ),
  .cpurst_b                             (cpurst_b                             ),
  .forever_cpuclk                       (forever_cpuclk                       ),
  .hpcp_cp0_cmplt                       (hpcp_cp0_cmplt                       ),
  .hpcp_cp0_data                        (hpcp_cp0_data                        ),
  .idu_cp0_rf_func                      (idu_cp0_rf_func                      ),
  .idu_cp0_rf_gateclk_sel               (idu_cp0_rf_gateclk_sel               ),
  .idu_cp0_rf_iid                       (idu_cp0_rf_iid                       ),
  .idu_cp0_rf_opcode                    (idu_cp0_rf_opcode                    ),
  .idu_cp0_rf_preg                      (idu_cp0_rf_preg                      ),
  .idu_cp0_rf_sel                       (idu_cp0_rf_sel                       ),
  .idu_cp0_rf_src0                      (idu_cp0_rf_src0                      ),
  .idu_cp0_rf_src1                      (idu_cp0_rf_src1                      ),
  .ifu_cp0_icache_inv_done              (ifu_cp0_icache_inv_done              ),
  .ifu_cp0_rst_inv_req                  (ifu_cp0_rst_inv_req                  ),
  .inst_lpmd_ex1_ex2                    (inst_lpmd_ex1_ex2                    ),
  .iui_regs_addr                        (iui_regs_addr                        ),
  .iui_regs_csr_wr                      (iui_regs_csr_wr                      ),
  .iui_regs_csrw                        (iui_regs_csrw                        ),
  .iui_regs_ex3_inst_csr                (iui_regs_ex3_inst_csr                ),
  .iui_regs_inst_mret                   (iui_regs_inst_mret                   ),
  .iui_regs_inst_ertn                   (iui_regs_inst_ertn                   ),
  .iui_regs_inst_sret                   (iui_regs_inst_sret                   ),
  .iui_regs_inv_expt                    (iui_regs_inv_expt                    ),
  .iui_regs_opcode                      (iui_regs_opcode                      ),
  .iui_regs_ori_src0                    (iui_regs_ori_src0                    ),
  .iui_regs_cpu_cfg_code                (iui_regs_cpu_cfg_code                ),
  .iui_regs_rst_inv_d                   (iui_regs_rst_inv_d                   ),
  .iui_regs_rst_inv_i                   (iui_regs_rst_inv_i                   ),
  .iui_regs_sel                         (iui_regs_sel                         ),
  .iui_regs_sel_ipi                     (iui_regs_sel_ipi                     ),
  .iui_regs_src0                        (iui_regs_src0                        ),
  .iui_regs_iocsr_addr                  (iui_regs_iocsr_addr                  ),
  .iui_ipi_regs_src                     (iui_ipi_regs_src                     ),
  .iui_update_ipi_status_en             (iui_update_ipi_status_en             ),
  .iui_update_ipi_status_src            (iui_update_ipi_status_src            ),
  .iui_update_ipi_mailbox0_en           (iui_update_ipi_mailbox0_en           ),
  .iui_update_ipi_mailbox1_en           (iui_update_ipi_mailbox1_en           ),
  .iui_update_ipi_mailbox2_en           (iui_update_ipi_mailbox2_en           ),
  .iui_update_ipi_mailbox3_en           (iui_update_ipi_mailbox3_en           ),
  .iui_update_ipi_mailbox_sel           (iui_update_ipi_mailbox_sel           ),
  .iui_update_ipi_regs_src0             (iui_update_ipi_regs_src0             ),
  .iui_update_ipi_regs_src1             (iui_update_ipi_regs_src1             ),
  .iui_update_ipi_regs_src2             (iui_update_ipi_regs_src2             ),
  .iui_update_ipi_regs_src3             (iui_update_ipi_regs_src3             ),
  .iui_update_ipi_regs_mask0            (iui_update_ipi_regs_mask0            ),
  .iui_update_ipi_regs_mask1            (iui_update_ipi_regs_mask1            ),
  .iui_update_ipi_regs_mask2            (iui_update_ipi_regs_mask2            ),
  .iui_update_ipi_regs_mask3            (iui_update_ipi_regs_mask3            ),
  .iui_top_cur_state                    (iui_top_cur_state                    ),
  .lpmd_cmplt                           (lpmd_cmplt                           ),
  .lsu_cp0_dcache_done                  (lsu_cp0_dcache_done                  ),
  .mmu_cp0_cmplt                        (mmu_cp0_cmplt                        ),
  .mmu_cp0_tlb_done                     (mmu_cp0_tlb_done                     ),
  .pad_yy_icg_scan_en                   (pad_yy_icg_scan_en                   ),
  .sysio_core_restart_vld               (sysio_core_restart_vld               ),
  .core_sysio_restart_grnt              (core_sysio_restart_grnt              ),
  .sysio_core_cp0_update_ipi_status_en  (sysio_core_cp0_update_ipi_status_en  ),
  .sysio_core_cp0_update_ipi_status_src (sysio_core_cp0_update_ipi_status_src ),
  .sysio_core_cp0_update_mailbox0_en    (sysio_core_cp0_update_mailbox0_en    ),
  .sysio_core_cp0_update_mailbox1_en    (sysio_core_cp0_update_mailbox1_en    ),
  .sysio_core_cp0_update_mailbox2_en    (sysio_core_cp0_update_mailbox2_en    ),
  .sysio_core_cp0_update_mailbox3_en    (sysio_core_cp0_update_mailbox3_en    ),
  .sysio_core_cp0_req_grnt              (sysio_core_cp0_req_grnt              ),
  .sysio_core_cp0_update_bit_sel        (sysio_core_cp0_update_bit_sel        ),
  .sysio_core_cp0_update_mailbox_src0   (sysio_core_cp0_update_mailbox_src0   ),
  .sysio_core_cp0_update_mailbox_src1   (sysio_core_cp0_update_mailbox_src1   ),
  .sysio_core_cp0_update_mailbox_src2   (sysio_core_cp0_update_mailbox_src2   ),
  .sysio_core_cp0_update_mailbox_src3   (sysio_core_cp0_update_mailbox_src3   ),
  .sysio_core_cp0_update_mailbox_mask0  (sysio_core_cp0_update_mailbox_mask0  ),
  .sysio_core_cp0_update_mailbox_mask1  (sysio_core_cp0_update_mailbox_mask1  ),
  .sysio_core_cp0_update_mailbox_mask2  (sysio_core_cp0_update_mailbox_mask2  ),
  .sysio_core_cp0_update_mailbox_mask3  (sysio_core_cp0_update_mailbox_mask3  ),
  .regs_iui_cfr_no_op                   (regs_iui_cfr_no_op                   ),
  .regs_iui_chk_vld                     (regs_iui_chk_vld                     ),
  .regs_iui_cindex_l2                   (regs_iui_cindex_l2                   ),
  .regs_iui_cins_no_op                  (regs_iui_cins_no_op                  ),
  .regs_iui_cskyee                      (regs_iui_cskyee                      ),
  .regs_iui_data_out                    (regs_iui_data_out                    ),
  .regs_iui_iocsr_data_out              (regs_iui_iocsr_data_out              ),
  .regs_iui_mailbox0_data               (regs_iui_mailbox0_data               ),
  .regs_iui_cfg_data_out                (regs_iui_cfg_data_out                ),
  .regs_iui_dca_sel                     (regs_iui_dca_sel                     ),
  .regs_iui_fs_off                      (regs_iui_fs_off                      ),
  .regs_iui_hpcp_regs_sel               (regs_iui_hpcp_regs_sel               ),
  .regs_iui_hpcp_scr_inv                (regs_iui_hpcp_scr_inv                ),
  .regs_iui_int_sel                     (regs_iui_int_sel                     ),
  .regs_iui_l2_regs_sel                 (regs_iui_l2_regs_sel                 ),
  .regs_iui_pm                          (regs_iui_pm                          ),
  .regs_iui_reg_idx                     (regs_iui_reg_idx                     ),
  .regs_iui_scnt_inv                    (regs_iui_scnt_inv                    ),
  .regs_iui_tee_ff                      (regs_iui_tee_ff                      ),
  .regs_iui_tee_vld                     (regs_iui_tee_vld                     ),
  .regs_iui_tsr                         (regs_iui_tsr                         ),
  .regs_iui_tvm                         (regs_iui_tvm                         ),
  .regs_iui_tw                          (regs_iui_tw                          ),
  .regs_iui_ucnt_inv                    (regs_iui_ucnt_inv                    ),
  .regs_iui_v                           (regs_iui_v                           ),
  .regs_iui_vs_off                      (regs_iui_vs_off                      ),
  .regs_iui_ecfg_vs                     (regs_iui_ecfg_vs                     ),
  .regs_iui_wdata                       (regs_iui_wdata                       ),
  .regs_xx_icg_en                       (regs_xx_icg_en                       ),
  .rtu_yy_xx_commit0                    (rtu_yy_xx_commit0                    ),
  .rtu_yy_xx_commit0_iid                (rtu_yy_xx_commit0_iid                ),
  .rtu_yy_xx_dbgon                      (rtu_yy_xx_dbgon                      ),
  .rtu_yy_xx_flush                      (rtu_yy_xx_flush                      )
);


// &Instance("ct_cp0_regs", "x_ct_cp0_regs"); @34
ct_cp0_regs  x_ct_cp0_regs (
  .biu_cp0_apb_base                (biu_cp0_apb_base               ),
  .biu_cp0_cmplt                   (biu_cp0_cmplt                  ),
  .biu_cp0_coreid                  (biu_cp0_coreid                 ),
  .ext_interrupt                   (ext_interrupt                  ),
  .biu_cp0_me_int                  (biu_cp0_me_int                 ),
  .biu_cp0_ms_int                  (biu_cp0_ms_int                 ),
  .biu_cp0_mt_int                  (biu_cp0_mt_int                 ),
  .biu_cp0_rdata                   (biu_cp0_rdata                  ),
  .biu_cp0_rvba                    (biu_cp0_rvba                   ),
  .biu_cp0_se_int                  (biu_cp0_se_int                 ),
  .biu_cp0_ss_int                  (biu_cp0_ss_int                 ),
  .biu_cp0_st_int                  (biu_cp0_st_int                 ),
  .cp0_biu_icg_en                  (cp0_biu_icg_en                 ),
  .cp0_had_cpuid_0                 (cp0_had_cpuid_0                ),
  .cp0_had_trace_pm_wdata          (cp0_had_trace_pm_wdata         ),
  .cp0_had_trace_pm_wen            (cp0_had_trace_pm_wen           ),
  .cp0_hpcp_icg_en                 (cp0_hpcp_icg_en                ),
  .cp0_hpcp_index                  (cp0_hpcp_index                 ),
  .cp0_hpcp_int_disable            (cp0_hpcp_int_disable           ),
  .cp0_hpcp_mcntwen                (cp0_hpcp_mcntwen               ),
  .cp0_hpcp_pmdm                   (cp0_hpcp_pmdm                  ),
  .cp0_hpcp_pmds                   (cp0_hpcp_pmds                  ),
  .cp0_hpcp_pmdu                   (cp0_hpcp_pmdu                  ),
  .cp0_hpcp_wdata                  (cp0_hpcp_wdata                 ),
  .cp0_idu_cskyee                  (cp0_idu_cskyee                 ),
  .cp0_idu_dlb_disable             (cp0_idu_dlb_disable            ),
  .cp0_idu_frm                     (cp0_idu_frm                    ),
  .cp0_idu_fs                      (cp0_idu_fs                     ),
  .cp0_idu_icg_en                  (cp0_idu_icg_en                 ),
  .cp0_idu_iq_bypass_disable       (cp0_idu_iq_bypass_disable      ),
  .cp0_idu_rob_fold_disable        (cp0_idu_rob_fold_disable       ),
  .cp0_idu_src2_fwd_disable        (cp0_idu_src2_fwd_disable       ),
  .cp0_idu_srcv2_fwd_disable       (cp0_idu_srcv2_fwd_disable      ),
  .cp0_idu_vill                    (cp0_idu_vill                   ),
  .cp0_idu_vs                      (cp0_idu_vs                     ),
  .cp0_idu_vstart                  (cp0_idu_vstart                 ),
  .cp0_idu_zero_delay_move_disable (cp0_idu_zero_delay_move_disable),
  .cp0_ifu_bht_en                  (cp0_ifu_bht_en                 ),
  .cp0_ifu_bht_inv                 (cp0_ifu_bht_inv                ),
  .cp0_ifu_btb_en                  (cp0_ifu_btb_en                 ),
  .cp0_ifu_btb_inv                 (cp0_ifu_btb_inv                ),
  .cp0_ifu_icache_en               (cp0_ifu_icache_en              ),
  .cp0_ifu_icache_inv              (cp0_ifu_icache_inv             ),
  .cp0_ifu_icache_pref_en          (cp0_ifu_icache_pref_en         ),
  .cp0_ifu_icache_read_index       (cp0_ifu_icache_read_index      ),
  .cp0_ifu_icache_read_req         (cp0_ifu_icache_read_req        ),
  .cp0_ifu_icache_read_tag         (cp0_ifu_icache_read_tag        ),
  .cp0_ifu_icache_read_way         (cp0_ifu_icache_read_way        ),
  .cp0_ifu_icg_en                  (cp0_ifu_icg_en                 ),
  .cp0_ifu_ind_btb_en              (cp0_ifu_ind_btb_en             ),
  .cp0_ifu_ind_btb_inv             (cp0_ifu_ind_btb_inv            ),
  .cp0_ifu_insde                   (cp0_ifu_insde                  ),
  .cp0_ifu_iwpe                    (cp0_ifu_iwpe                   ),
  .cp0_ifu_l0btb_en                (cp0_ifu_l0btb_en               ),
  .cp0_ifu_lbuf_en                 (cp0_ifu_lbuf_en                ),
  .cp0_ifu_nsfe                    (cp0_ifu_nsfe                   ),
  .cp0_ifu_ras_en                  (cp0_ifu_ras_en                 ),
  .cp0_ifu_rvbr                    (cp0_ifu_rvbr                   ),
  .cp0_ifu_vbr                     (cp0_ifu_vbr                    ),
  .cp0_ifu_ecfg_vs                 (cp0_ifu_ecfg_vs                ),
  .cp0_ifu_eentry                  (cp0_ifu_eentry                 ),
  .cp0_ifu_vl                      (cp0_ifu_vl                     ),
  .cp0_ifu_vlmul                   (cp0_ifu_vlmul                  ),
  .cp0_ifu_vsetvli_pred_disable    (cp0_ifu_vsetvli_pred_disable   ),
  .cp0_ifu_vsetvli_pred_mode       (cp0_ifu_vsetvli_pred_mode      ),
  .cp0_ifu_vsew                    (cp0_ifu_vsew                   ),
  .cp0_iu_div_entry_disable        (cp0_iu_div_entry_disable       ),
  .cp0_iu_div_entry_disable_clr    (cp0_iu_div_entry_disable_clr   ),
  .cp0_iu_ex3_efpc                 (cp0_iu_ex3_efpc                ),
  .cp0_iu_ex3_efpc_vld             (cp0_iu_ex3_efpc_vld            ),
  .cp0_iu_icg_en                   (cp0_iu_icg_en                  ),
  .cp0_iu_bju_chflw_en             (cp0_iu_bju_chflw_en            ),
  .cp0_iu_vill                     (cp0_iu_vill                    ),
  .cp0_iu_vl                       (cp0_iu_vl                      ),
  .cp0_iu_vsetvli_pre_decd_disable (cp0_iu_vsetvli_pre_decd_disable),
  .cp0_iu_vstart                   (cp0_iu_vstart                  ),
  .cp0_iu_timer                    (cp0_iu_timer                   ),
  .cp0_lsu_amr                     (cp0_lsu_amr                    ),
  .cp0_lsu_amr2                    (cp0_lsu_amr2                   ),
  .cp0_lsu_cb_aclr_dis             (cp0_lsu_cb_aclr_dis            ),
  .cp0_lsu_corr_dis                (cp0_lsu_corr_dis               ),
  .cp0_lsu_ctc_flush_dis           (cp0_lsu_ctc_flush_dis          ),
  .cp0_lsu_da_fwd_dis              (cp0_lsu_da_fwd_dis             ),
  .cp0_lsu_dcache_clr              (cp0_lsu_dcache_clr             ),
  .cp0_lsu_dcache_en               (cp0_lsu_dcache_en              ),
  .cp0_lsu_dcache_inv              (cp0_lsu_dcache_inv             ),
  .cp0_lsu_dcache_pref_dist        (cp0_lsu_dcache_pref_dist       ),
  .cp0_lsu_dcache_pref_en          (cp0_lsu_dcache_pref_en         ),
  .cp0_lsu_dcache_read_index       (cp0_lsu_dcache_read_index      ),
  .cp0_lsu_dcache_read_ld_tag      (cp0_lsu_dcache_read_ld_tag     ),
  .cp0_lsu_dcache_read_req         (cp0_lsu_dcache_read_req        ),
  .cp0_lsu_dcache_read_st_tag      (cp0_lsu_dcache_read_st_tag     ),
  .cp0_lsu_dcache_read_way         (cp0_lsu_dcache_read_way        ),
  .cp0_lsu_fencei_broad_dis        (cp0_lsu_fencei_broad_dis       ),
  .cp0_lsu_fencerw_broad_dis       (cp0_lsu_fencerw_broad_dis      ),
  .cp0_lsu_icg_en                  (cp0_lsu_icg_en                 ),
  .cp0_lsu_l2_pref_dist            (cp0_lsu_l2_pref_dist           ),
  .cp0_lsu_l2_pref_en              (cp0_lsu_l2_pref_en             ),
  .cp0_lsu_l2_st_pref_en           (cp0_lsu_l2_st_pref_en          ),
  .cp0_lsu_mm                      (cp0_lsu_mm                     ),
  .cp0_lsu_nsfe                    (cp0_lsu_nsfe                   ),
  .cp0_lsu_pfu_mmu_dis             (cp0_lsu_pfu_mmu_dis            ),
  .cp0_lsu_timeout_cnt             (cp0_lsu_timeout_cnt            ),
  .cp0_lsu_tlb_broad_dis           (cp0_lsu_tlb_broad_dis          ),
  .cp0_lsu_tvm                     (cp0_lsu_tvm                    ),
  .cp0_lsu_ucme                    (cp0_lsu_ucme                   ),
  .cp0_lsu_vstart                  (cp0_lsu_vstart                 ),
  .cp0_lsu_wa                      (cp0_lsu_wa                     ),
  .cp0_lsu_wr_burst_dis            (cp0_lsu_wr_burst_dis           ),
  .cp0_mmu_cskyee                  (cp0_mmu_cskyee                 ),
  .cp0_mmu_icg_en                  (cp0_mmu_icg_en                 ),
  .cp0_mmu_maee                    (cp0_mmu_maee                   ),
  .cp0_mmu_mpp                     (cp0_mmu_mpp                    ),
  .cp0_mmu_mprv                    (cp0_mmu_mprv                   ),
  .cp0_mmu_mxr                     (cp0_mmu_mxr                    ),
  .cp0_mmu_ptw_en                  (cp0_mmu_ptw_en                 ),
  .cp0_mmu_reg_num                 (cp0_mmu_reg_num                ),
  .cp0_mmu_satp_sel                (cp0_mmu_satp_sel               ),
  .cp0_mmu_sum                     (cp0_mmu_sum                    ),
  .cp0_mmu_wdata                   (cp0_mmu_wdata                  ),
  .cp0_mmu_wreg                    (cp0_mmu_wreg                   ),
  .cp0_mmu_crmd_da                 (cp0_mmu_crmd_da                ),
  .cp0_mmu_crmd_pg                 (cp0_mmu_crmd_pg                ),
  .cp0_mmu_cur_asid                (cp0_mmu_cur_asid               ),
  .cp0_mmu_da_mode_datf            (cp0_mmu_da_mode_datf           ),
  .cp0_mmu_da_mode_datm            (cp0_mmu_da_mode_datm           ),
  .cp0_mmu_ptw_pgdl                (cp0_mmu_ptw_pgdl               ),
  .cp0_mmu_ptw_pgdh                (cp0_mmu_ptw_pgdh               ),
  .cp0_mmu_dmw0                    (cp0_mmu_dmw0                   ),
  .cp0_mmu_dmw1                    (cp0_mmu_dmw1                   ),
  .cp0_mmu_dmw2                    (cp0_mmu_dmw2                   ),
  .cp0_mmu_dmw3                    (cp0_mmu_dmw3                   ),
  .cp0_mret                        (cp0_mret                       ),
  .cp0_ertn                        (cp0_ertn                       ),
  .cp0_cprs                        (cp0_cprs                       ),
  .cp0_pad_mstatus                 (cp0_pad_mstatus                ),
  .cp0_pmp_icg_en                  (cp0_pmp_icg_en                 ),
  .cp0_pmp_mpp                     (cp0_pmp_mpp                    ),
  .cp0_pmp_mprv                    (cp0_pmp_mprv                   ),
  .cp0_pmp_reg_num                 (cp0_pmp_reg_num                ),
  .cp0_pmp_wdata                   (cp0_pmp_wdata                  ),
  .cp0_pmp_wreg                    (cp0_pmp_wreg                   ),
  .cp0_rtu_icg_en                  (cp0_rtu_icg_en                 ),
  .cp0_rtu_srt_en                  (cp0_rtu_srt_en                 ),
  .cp0_sret                        (cp0_sret                       ),
  .cp0_vfpu_fcsr                   (cp0_vfpu_fcsr                  ),
  .cp0_vfpu_fxcr                   (cp0_vfpu_fxcr                  ),
  .cp0_vfpu_icg_en                 (cp0_vfpu_icg_en                ),
  .cp0_vfpu_vl                     (cp0_vfpu_vl                    ),
  .cp0_xx_core_arch                (cp0_xx_core_arch               ),
  .cp0_xx_core_icg_en              (cp0_xx_core_icg_en             ),
  .cp0_yy_clk_en                   (cp0_yy_clk_en                  ),
  .cp0_yy_dcache_pref_en           (cp0_yy_dcache_pref_en          ),
  .cp0_yy_hyper                    (cp0_yy_hyper                   ),
  .cp0_yy_priv_mode                (cp0_yy_priv_mode               ),
  .cp0_yy_virtual_mode             (cp0_yy_virtual_mode            ),
  .cpurst_b                        (cpurst_b                       ),
  .forever_cpuclk                  (forever_cpuclk                 ),
  .hpcp_cp0_data                   (hpcp_cp0_data                  ),
  .hpcp_cp0_int_vld                (hpcp_cp0_int_vld               ),
  .hpcp_cp0_sce                    (hpcp_cp0_sce                   ),
  .idu_cp0_fesr_acc_updt_val       (idu_cp0_fesr_acc_updt_val      ),
  .idu_cp0_fesr_acc_updt_vld       (idu_cp0_fesr_acc_updt_vld      ),
  .ifu_cp0_bht_inv_done            (ifu_cp0_bht_inv_done           ),
  .ifu_cp0_btb_inv_done            (ifu_cp0_btb_inv_done           ),
  .ifu_cp0_icache_inv_done         (ifu_cp0_icache_inv_done        ),
  .ifu_cp0_icache_read_data        (ifu_cp0_icache_read_data       ),
  .ifu_cp0_icache_read_data_vld    (ifu_cp0_icache_read_data_vld   ),
  .ifu_cp0_ind_btb_inv_done        (ifu_cp0_ind_btb_inv_done       ),
  .ifu_cp0_rst_inv_req             (ifu_cp0_rst_inv_req            ),
  .iui_regs_addr                   (iui_regs_addr                  ),
  .iui_regs_csr_wr                 (iui_regs_csr_wr                ),
  .iui_regs_csrw                   (iui_regs_csrw                  ),
  .iui_regs_ex3_inst_csr           (iui_regs_ex3_inst_csr          ),
  .iui_regs_inst_mret              (iui_regs_inst_mret             ),
  .iui_regs_inst_ertn              (iui_regs_inst_ertn             ),
  .iui_regs_inst_sret              (iui_regs_inst_sret             ),
  .iui_regs_inv_expt               (iui_regs_inv_expt              ),
  .iui_regs_opcode                 (iui_regs_opcode                ),
  .iui_regs_ori_src0               (iui_regs_ori_src0              ),
  .iui_regs_cpu_cfg_code           (iui_regs_cpu_cfg_code          ),
  .iui_regs_rst_inv_d              (iui_regs_rst_inv_d             ),
  .iui_regs_rst_inv_i              (iui_regs_rst_inv_i             ),
  .iui_regs_sel                    (iui_regs_sel                   ),
  .iui_regs_sel_ipi                (iui_regs_sel_ipi               ),
  .iui_regs_src0                   (iui_regs_src0                  ),
  .iui_ipi_regs_src                (iui_ipi_regs_src               ),
  .iui_regs_iocsr_addr             (iui_regs_iocsr_addr            ),
  .iui_update_ipi_status_en        (iui_update_ipi_status_en       ),
  .iui_update_ipi_status_src       (iui_update_ipi_status_src      ),
  .iui_update_ipi_mailbox0_en      (iui_update_ipi_mailbox0_en     ),
  .iui_update_ipi_mailbox1_en      (iui_update_ipi_mailbox1_en     ),
  .iui_update_ipi_mailbox2_en      (iui_update_ipi_mailbox2_en     ),
  .iui_update_ipi_mailbox3_en      (iui_update_ipi_mailbox3_en     ),
  .iui_update_ipi_mailbox_sel      (iui_update_ipi_mailbox_sel     ),
  .iui_update_ipi_regs_src0        (iui_update_ipi_regs_src0       ),
  .iui_update_ipi_regs_src1        (iui_update_ipi_regs_src1       ),
  .iui_update_ipi_regs_src2        (iui_update_ipi_regs_src2       ),
  .iui_update_ipi_regs_src3        (iui_update_ipi_regs_src3       ),
  .iui_update_ipi_regs_mask0       (iui_update_ipi_regs_mask0      ),
  .iui_update_ipi_regs_mask1       (iui_update_ipi_regs_mask1      ),
  .iui_update_ipi_regs_mask2       (iui_update_ipi_regs_mask2      ),
  .iui_update_ipi_regs_mask3       (iui_update_ipi_regs_mask3      ),
  .lsu_cp0_dcache_done             (lsu_cp0_dcache_done            ),
  .lsu_cp0_dcache_read_data        (lsu_cp0_dcache_read_data       ),
  .lsu_cp0_dcache_read_data_vld    (lsu_cp0_dcache_read_data_vld   ),
  .lsu_cp0_ld_va                   (lsu_cp0_ld_va                  ),
  .lsu_cp0_ld_pa                   (lsu_cp0_ld_pa                  ),
  .lsu_cp0_ld_vld                  (lsu_cp0_ld_vld                 ),
  .mmu_cp0_data                    (mmu_cp0_data                   ),
  .mmu_cp0_satp_data               (mmu_cp0_satp_data              ),
  .mmu_cp0_type                    (mmu_cp0_type                   ),
  .mmu_cp0_vpn                     (mmu_cp0_vpn                    ),
  .mmu_cp0_fst_vld                 (mmu_cp0_fst_vld                ),
  .mmu_cp0_fst_addr                (mmu_cp0_fst_addr               ),
  .mmu_cp0_scd_vld                 (mmu_cp0_scd_vld                ),
  .mmu_cp0_scd_addr                (mmu_cp0_scd_addr               ),
  .mmu_cp0_thd_vld                 (mmu_cp0_thd_vld                ),
  .mmu_cp0_thd_addr                (mmu_cp0_thd_addr               ),
  .pad_yy_icg_scan_en              (pad_yy_icg_scan_en             ),
  .pmp_cp0_data                    (pmp_cp0_data                   ),
  .sysio_core_gl_stable_timer      (sysio_core_gl_stable_timer     ),
  .regs_iui_cfr_no_op              (regs_iui_cfr_no_op             ),
  .regs_iui_chk_vld                (regs_iui_chk_vld               ),
  .regs_iui_cindex_l2              (regs_iui_cindex_l2             ),
  .regs_iui_cins_no_op             (regs_iui_cins_no_op            ),
  .regs_iui_cskyee                 (regs_iui_cskyee                ),
  .regs_iui_data_out               (regs_iui_data_out              ),
  .regs_iui_iocsr_data_out         (regs_iui_iocsr_data_out        ),
  .regs_iui_mailbox0_data          (regs_iui_mailbox0_data         ),
  .regs_iui_cfg_data_out           (regs_iui_cfg_data_out          ),
  .regs_iui_dca_sel                (regs_iui_dca_sel               ),
  .regs_iui_fs_off                 (regs_iui_fs_off                ),
  .regs_iui_hpcp_regs_sel          (regs_iui_hpcp_regs_sel         ),
  .regs_iui_hpcp_scr_inv           (regs_iui_hpcp_scr_inv          ),
  .regs_iui_int_sel                (regs_iui_int_sel               ),
  .regs_iui_l2_regs_sel            (regs_iui_l2_regs_sel           ),
  .regs_iui_pm                     (regs_iui_pm                    ),
  .regs_iui_reg_idx                (regs_iui_reg_idx               ),
  .regs_iui_scnt_inv               (regs_iui_scnt_inv              ),
  .regs_iui_tee_ff                 (regs_iui_tee_ff                ),
  .regs_iui_tee_vld                (regs_iui_tee_vld               ),
  .regs_iui_tsr                    (regs_iui_tsr                   ),
  .regs_iui_tvm                    (regs_iui_tvm                   ),
  .regs_iui_tw                     (regs_iui_tw                    ),
  .regs_iui_ucnt_inv               (regs_iui_ucnt_inv              ),
  .regs_iui_v                      (regs_iui_v                     ),
  .regs_iui_vs_off                 (regs_iui_vs_off                ),
  .regs_iui_ecfg_vs                (regs_iui_ecfg_vs               ),
  .regs_iui_wdata                  (regs_iui_wdata                 ),
  .regs_lpmd_int_vld               (regs_lpmd_int_vld              ),
  .regs_xx_icg_en                  (regs_xx_icg_en                 ),
  .rtu_cp0_epc                     (rtu_cp0_epc                    ),
  .rtu_cp0_expt_gateclk_vld        (rtu_cp0_expt_gateclk_vld       ),
  .rtu_cp0_expt_mtval              (rtu_cp0_expt_mtval             ),
  .rtu_cp0_expt_vld                (rtu_cp0_expt_vld               ),
  .rtu_cp0_fp_dirty_vld            (rtu_cp0_fp_dirty_vld           ),
  .rtu_cp0_int_ack                 (rtu_cp0_int_ack                ),
  .rtu_cp0_vec_dirty_vld           (rtu_cp0_vec_dirty_vld          ),
  .rtu_cp0_vsetvl_vill             (rtu_cp0_vsetvl_vill            ),
  .rtu_cp0_vsetvl_vl               (rtu_cp0_vsetvl_vl              ),
  .rtu_cp0_vsetvl_vl_vld           (rtu_cp0_vsetvl_vl_vld          ),
  .rtu_cp0_vsetvl_vlmul            (rtu_cp0_vsetvl_vlmul           ),
  .rtu_cp0_vsetvl_vsew             (rtu_cp0_vsetvl_vsew            ),
  .rtu_cp0_vsetvl_vtype_vld        (rtu_cp0_vsetvl_vtype_vld       ),
  .rtu_cp0_vstart                  (rtu_cp0_vstart                 ),
  .rtu_cp0_vstart_vld              (rtu_cp0_vstart_vld             ),
  .rtu_yy_xx_expt_vec              (rtu_yy_xx_expt_vec             ),
  .rtu_yy_xx_flush                 (rtu_yy_xx_flush                )
);


// &Instance("ct_cp0_lpmd", "x_ct_cp0_lpmd"); @36
ct_cp0_lpmd  x_ct_cp0_lpmd (
  .biu_yy_xx_no_op    (biu_yy_xx_no_op   ),
  .cp0_biu_lpmd_b     (cp0_biu_lpmd_b    ),
  .cp0_had_lpmd_b     (cp0_had_lpmd_b    ),
  .cp0_ifu_no_op_req  (cp0_ifu_no_op_req ),
  .cp0_lsu_no_op_req  (cp0_lsu_no_op_req ),
  .cp0_mmu_no_op_req  (cp0_mmu_no_op_req ),
  .cp0_yy_clk_en      (cp0_yy_clk_en     ),
  .cpurst_b           (cpurst_b          ),
  .forever_cpuclk     (forever_cpuclk    ),
  .had_cp0_xx_dbg     (had_cp0_xx_dbg    ),
  .ifu_yy_xx_no_op    (ifu_yy_xx_no_op   ),
  .inst_lpmd_ex1_ex2  (inst_lpmd_ex1_ex2 ),
  .lpmd_cmplt         (lpmd_cmplt        ),
  .lpmd_top_cur_state (lpmd_top_cur_state),
  .lsu_yy_xx_no_op    (lsu_yy_xx_no_op   ),
  .mmu_yy_xx_no_op    (mmu_yy_xx_no_op   ),
  .pad_yy_icg_scan_en (pad_yy_icg_scan_en),
  .regs_lpmd_int_vld  (regs_lpmd_int_vld ),
  .regs_xx_icg_en     (regs_xx_icg_en    ),
  .rtu_yy_xx_dbgon    (rtu_yy_xx_dbgon   ),
  .rtu_yy_xx_flush    (rtu_yy_xx_flush   )
);


assign cp0_had_debug_info[1:0] = iui_top_cur_state[1:0];
assign cp0_had_debug_info[3:2] = lpmd_top_cur_state[1:0];

// //&Force("nonport","mp_lpmd"); @143
// //&Force("nonport","mp_rst_b"); @144
// //&Force("nonport","mp_wakeup"); @145

// &ModuleEnd; @178
endmodule



