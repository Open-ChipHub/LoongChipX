`timescale 1ns/1ps 

module Sim_Top #(
    parameter int unsigned AXI_ID_WIDTH      = 8,
    parameter int unsigned AXI_ADDR_WIDTH    = 40,
    parameter int unsigned AXI_DATA_WIDTH    = 128,
    parameter int unsigned AXI_USER_WIDTH    = 2
)(
  output   wire                          axi_ar_valid,
  input    wire                          axi_ar_ready,
  output   wire   [AXI_ADDR_WIDTH-1:0]   axi_ar_addr,
  output   wire   [AXI_ID_WIDTH-1  :0]   axi_ar_id,
  output   wire   [7:0]                  axi_ar_len,
  output   wire   [2:0]                  axi_ar_size,
  output   wire   [1:0]                  axi_ar_burst,
  output   wire   [3:0]                  axi_ar_cache,
  output   wire   [2:0]                  axi_ar_prot,
  output   wire                          axi_aw_valid,
  input    wire                          axi_aw_ready,
  output   wire   [AXI_ADDR_WIDTH-1:0]   axi_aw_addr,
  output   wire   [AXI_ID_WIDTH-1  :0]   axi_aw_id,
  output   wire   [7:0]                  axi_aw_len,
  output   wire   [2:0]                  axi_aw_size,
  output   wire   [1:0]                  axi_aw_burst,
  output   wire   [3:0]                  axi_aw_cache,
  output   wire   [2:0]                  axi_aw_prot,
  output   wire                          axi_w_valid,
  input    wire                          axi_w_ready,
  output   wire   [AXI_DATA_WIDTH-1:0]   axi_w_data,
  output   wire   [15:0]                 axi_w_strb,
  output   wire                          axi_w_last,
  input    wire                          axi_b_valid,
  output   wire                          axi_b_ready,
  input    wire   [AXI_ID_WIDTH-1  :0]   axi_b_id,
  input    wire   [1:0]                  axi_b_resp,
  input    wire                          axi_r_valid,
  output   wire                          axi_r_ready,
  input    wire   [AXI_DATA_WIDTH-1:0]   axi_r_data,
  input    wire   [AXI_ID_WIDTH-1  :0]   axi_r_id,
  input    wire   [1:0]                  axi_r_resp,
  input    wire                          axi_r_last,
  input    wire   [7:0]                  core_in_interrupt,
  input    wire                          reset,
  input    wire                          clk
);

Top Top (
  .axi_ar_valid (axi_ar_valid),
  .axi_ar_ready (axi_ar_ready),
  .axi_ar_addr  (axi_ar_addr),
  .axi_ar_id    (axi_ar_id),
  .axi_ar_len   (axi_ar_len),
  .axi_ar_size  (axi_ar_size),
  .axi_ar_burst (axi_ar_burst),
  .axi_ar_cache (axi_ar_cache),
  .axi_ar_prot  (axi_ar_prot),
  .axi_aw_valid (axi_aw_valid),
  .axi_aw_ready (axi_aw_ready),
  .axi_aw_addr  (axi_aw_addr),
  .axi_aw_id    (axi_aw_id),
  .axi_aw_len   (axi_aw_len),
  .axi_aw_size  (axi_aw_size),
  .axi_aw_burst (axi_aw_burst),
  .axi_aw_cache (axi_aw_cache),
  .axi_aw_prot  (axi_aw_prot),
  .axi_w_valid  (axi_w_valid),
  .axi_w_ready  (axi_w_ready),
  .axi_w_data   (axi_w_data),
  .axi_w_strb   (axi_w_strb),
  .axi_w_last   (axi_w_last),
  .axi_b_valid  (axi_b_valid),
  .axi_b_ready  (axi_b_ready),
  .axi_b_id     (axi_b_id),
  .axi_b_resp   (axi_b_resp),
  .axi_r_valid  (axi_r_valid),
  .axi_r_ready  (axi_r_ready),
  .axi_r_data   (axi_r_data),
  .axi_r_id     (axi_r_id),
  .axi_r_resp   (axi_r_resp),
  .axi_r_last   (axi_r_last),
  .core_in_interrupt (core_in_interrupt),
  .dbg_sim_cycles(),
  .reset        (reset),
  .clk          (clk)
  );

endmodule