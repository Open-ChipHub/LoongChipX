/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @23
module aq_ifu_pcgen (
  // &Ports, @24
  input    wire  [63:0]  btb_pcgen_tar_pc,
  input    wire          btb_xx_chgflw_vld,
  input    wire          cp0_ifu_icg_en,
  input    wire  [63:0]  cp0_xx_mrvbr,
  input    wire          cp0_yy_clk_en,
  input    wire          cpurst_b,
  input    wire          forever_cpuclk,
  input    wire  [63:0]  icache_pcgen_addr,
  input    wire          icache_pcgen_grant,
  input    wire          icache_pcgen_grant_gate,
  input    wire          icache_pcgen_inst_vld,
  input    wire          icache_pcgen_inst_vld_gate,
  input    wire          ipack_pcgen_reissue,
  input    wire  [63:0]  iu_ifu_tar_pc,
  input    wire          iu_ifu_tar_pc_vld,
  input    wire          iu_ifu_tar_pc_vld_gate,
  input    wire          pad_yy_icg_scan_en,
  input    wire  [63:0]  pred_pcgen_chgflw_pc,
  input    wire          pred_pcgen_chgflw_vld,
  input    wire          pred_pcgen_chgflw_vld_gate,
  input    wire  [63:0]  pred_pcgen_curflw_pc,
  input    wire          pred_pcgen_curflw_vld,
  input    wire          pred_pcgen_curflw_vld_gate,
  input    wire  [63:0]  rtu_ifu_chgflw_pc,
  input    wire          rtu_ifu_chgflw_vld,
  input    wire          vec_pcgen_idle,
  input    wire          vec_pcgen_rst_vld,
  output   wire  [63:0]  ifu_iu_chgflw_pc,
  output   wire          ifu_iu_chgflw_vld,
  output   wire  [63:0]  pcgen_btb_ifpc,
  output   wire          pcgen_ctrl_chgflw_vld,
  output   wire          pcgen_ibuf_chgflw_vld,
  output   wire          pcgen_icache_chgflw_vld,
  output   wire  [33:0]  pcgen_icache_seq_tag,
  output   wire  [63:0]  pcgen_icache_va,
  output   wire          pcgen_pred_flush_vld,
  output   wire  [63:0]  pcgen_pred_ifpc,
  output   wire          pcgen_top_buf_chgflw
); 



// &Regs; @25
reg             pcgen_buf_chgflw;           
reg     [63:0]  pcgen_ifpc;                 
reg     [63:0]  pcgen_pipe_ifpc;            

// &Wires; @26
wire    [63:0]  pcgen_br_chgflw_pc;         
wire            pcgen_br_chgflw_vld;        
wire            pcgen_chgflw_btb;           
wire            pcgen_chgflw_cur;           
wire            pcgen_cpuclk;               
wire    [63:0]  pcgen_delay_chgflw_pc;      
wire            pcgen_delay_chgflw_vld;     
wire            pcgen_delay_chgflw_vld_gate; 
wire    [63:0]  pcgen_fetch_pc;             
wire            pcgen_icg_en;               
wire    [63:0]  pcgen_ifpc_inc;             


//==========================================================
// PC Generator Module
// 1. ICG Instance
// 2. Judge the priority of PC sources
// 3. IF PC Maintain
//==========================================================

//------------------------------------------------
// 1. ICG Instance
//------------------------------------------------
assign pcgen_icg_en = pcgen_delay_chgflw_vld_gate
                   || pcgen_buf_chgflw
                   || pred_pcgen_curflw_vld_gate
                   || btb_xx_chgflw_vld
                   || icache_pcgen_inst_vld_gate
                   || icache_pcgen_grant_gate
                   || vec_pcgen_rst_vld;
// &Instance("gated_clk_cell", "x_ifu_pcgen_icg_cell"); @45
gated_clk_cell  x_ifu_pcgen_icg_cell (
  .clk_in             (forever_cpuclk    ),
  .clk_out            (pcgen_cpuclk      ),
  .external_en        (1'b0              ),
  .global_en          (cp0_yy_clk_en     ),
  .local_en           (pcgen_icg_en      ),
  .module_en          (cp0_ifu_icg_en    ),
  .pad_yy_icg_scan_en (pad_yy_icg_scan_en)
);

// &Connect(.clk_in      (forever_cpuclk), @46
//          .external_en (1'b0), @47
//          .global_en   (cp0_yy_clk_en), @48
//          .module_en   (cp0_ifu_icg_en), @49
//          .local_en    (pcgen_icg_en), @50
//          .clk_out     (pcgen_cpuclk) @51
//        ); @52

//assign pcgen_high_icg_en = iu_ifu_tar_pc_vld
//                        || pcgen_high_upd
//                        || vec_pcgen_rst_vld;
//&Instance("gated_clk_cell", "x_ifu_pcgen_high_icg_cell");
// //&Connect(.clk_in      (forever_cpuclk), @58
// //         .external_en (1'b0), @59
// //         .global_en   (cp0_yy_clk_en), @60
// //         .module_en   (1'b0), @61
// //         .local_en    (pcgen_high_icg_en), @62
// //         .clk_out     (pcgen_high_cpuclk) @63
// //       ); @64
//------------------------------------------------
// 2. Judge the priority of PC sources
// a. Delayed change flow: RTU > BJU > Pred
// b. Normal change flow: BTB > Inc
//------------------------------------------------
// a. Delayed change flow: RTU > BJU > Pred
// Following change flow are delayed for timing
assign pcgen_br_chgflw_vld      = (iu_ifu_tar_pc_vld || pred_pcgen_chgflw_vld)
                               && !rtu_ifu_chgflw_vld;
assign pcgen_br_chgflw_pc[63:0] = iu_ifu_tar_pc_vld ? iu_ifu_tar_pc[63:0]
                                                    : pred_pcgen_chgflw_pc[63:0];
assign pcgen_delay_chgflw_vld      = rtu_ifu_chgflw_vld
                                  || iu_ifu_tar_pc_vld
                                  || pred_pcgen_chgflw_vld;
assign pcgen_delay_chgflw_vld_gate = rtu_ifu_chgflw_vld
                                  || iu_ifu_tar_pc_vld_gate
                                  || pred_pcgen_chgflw_vld_gate;
assign pcgen_delay_chgflw_pc[63:0] = {64{rtu_ifu_chgflw_vld}}  & rtu_ifu_chgflw_pc[63:0]
                                   | {64{pcgen_br_chgflw_vld}} & pcgen_br_chgflw_pc[63:0];

always @ (posedge pcgen_cpuclk or negedge cpurst_b)
begin
  if(!cpurst_b)
    pcgen_buf_chgflw <= 1'b0;
  else if(pcgen_delay_chgflw_vld)
    pcgen_buf_chgflw <= 1'b1;
  else if(pcgen_buf_chgflw)
    pcgen_buf_chgflw <= 1'b0;
end

//------------------------------------------------
// 3. IF PC Maintain
// a. Normal IFPC for 40-bit Virtual PC
// b. High IFPC for 64-bit PC validation
//------------------------------------------------
// a. Normal IFPC for 40-bit Virtual PC
always @ (posedge pcgen_cpuclk)
begin
  if(vec_pcgen_rst_vld)
    pcgen_ifpc[63:0] <= cp0_xx_mrvbr[63:0];
  else if(pcgen_delay_chgflw_vld)
    pcgen_ifpc[63:0] <= pcgen_delay_chgflw_pc[63:0];
  else if(pcgen_chgflw_cur && !icache_pcgen_grant)
    pcgen_ifpc[63:0] <= pcgen_fetch_pc[63:0];
  else if(ipack_pcgen_reissue && icache_pcgen_inst_vld)
    pcgen_ifpc[63:0] <= icache_pcgen_addr[63:0];
  else if(pcgen_chgflw_btb && !icache_pcgen_grant)
    pcgen_ifpc[63:0] <= pcgen_fetch_pc[63:0];
  else if(icache_pcgen_grant)
    pcgen_ifpc[63:0] <= pcgen_ifpc_inc[63:0];
  else
    pcgen_ifpc[63:0] <= pcgen_ifpc[63:0];
end

assign pcgen_ifpc_inc[63:0] = {pcgen_fetch_pc[63:2], 2'b0} + 64'h4;

assign pcgen_chgflw_btb     = btb_xx_chgflw_vld && !pcgen_buf_chgflw;
assign pcgen_chgflw_cur     = pred_pcgen_curflw_vld && !pcgen_buf_chgflw;
assign pcgen_fetch_pc[63:0] = pcgen_chgflw_cur ? {pred_pcgen_curflw_pc[63:0]}
                            : pcgen_chgflw_btb ? {btb_pcgen_tar_pc[63:0]}
                                               : pcgen_ifpc[63:0];

always @ (posedge pcgen_cpuclk)
begin
  if(vec_pcgen_rst_vld)
    pcgen_pipe_ifpc[63:0] <= cp0_xx_mrvbr[63:0];
  else if(icache_pcgen_grant)
    pcgen_pipe_ifpc[63:0] <= pcgen_fetch_pc[63:0];
  else
    pcgen_pipe_ifpc[63:0] <= pcgen_pipe_ifpc[63:0];
end

//==========================================================
// Rename for Output
//==========================================================

// Output to Ctrl
assign pcgen_ctrl_chgflw_vld = pcgen_delay_chgflw_vld || pred_pcgen_curflw_vld
                            || pcgen_buf_chgflw;

// Output to I-Buf
assign pcgen_ibuf_chgflw_vld = rtu_ifu_chgflw_vld
                            || iu_ifu_tar_pc_vld;

// Output to ICACHE
assign pcgen_icache_chgflw_vld = pcgen_delay_chgflw_vld || pred_pcgen_curflw_vld
                              || pcgen_buf_chgflw || btb_xx_chgflw_vld;
assign pcgen_icache_va[63:0]   = pcgen_fetch_pc[63:0];
assign pcgen_icache_seq_tag[33:0] = pcgen_ifpc[39:6];

// Output to BTB
assign pcgen_btb_ifpc[63:0]  = {pcgen_ifpc[63:16], pcgen_fetch_pc[15:0]};

// Output to Prediction
assign pcgen_pred_flush_vld  = rtu_ifu_chgflw_vld
                            || iu_ifu_tar_pc_vld;
assign pcgen_pred_ifpc[63:0] = pcgen_pipe_ifpc[63:0];

// Output to Top
assign pcgen_top_buf_chgflw  = pcgen_buf_chgflw;

// Output to IU
assign ifu_iu_chgflw_vld      = rtu_ifu_chgflw_vld;
assign ifu_iu_chgflw_pc[63:0] = pcgen_delay_chgflw_pc[63:0];

// &Force("input", "vec_pcgen_idle"); @192
// &Force("nonport", "rst_done"); @194

// &ModuleEnd; @224
endmodule


