/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @23
module aq_rtu_top (
  // &Ports, @25
  input    wire          cp0_rtu_ex1_chgflw,
  input    wire  [63:0]  cp0_rtu_ex1_chgflw_pc,
  input    wire          cp0_rtu_ex1_cmplt,
  input    wire          cp0_rtu_ex1_cmplt_dp,
  input    wire  [63:0]  cp0_rtu_ex1_expt_tval,
  input    wire  [14:0]  cp0_rtu_ex1_expt_vec,
  input    wire          cp0_rtu_ex1_expt_vld,
  input    wire          cp0_rtu_ex1_flush,
  input    wire  [21:0]  cp0_rtu_ex1_halt_info,
  input    wire          cp0_rtu_ex1_inst_dret,
  input    wire          cp0_rtu_ex1_inst_ebreak,
  input    wire          cp0_rtu_ex1_inst_len,
  input    wire          cp0_rtu_ex1_inst_ertn,
  input    wire          cp0_rtu_ex1_inst_mret,
  input    wire          cp0_rtu_ex1_inst_split,
  input    wire          cp0_rtu_ex1_inst_sret,
  input    wire          cp0_rtu_ex1_vs_dirty,
  input    wire          cp0_rtu_ex1_vs_dirty_dp,
  input    wire  [63:0]  cp0_rtu_ex1_wb_data,
  input    wire          cp0_rtu_ex1_wb_dp,
  input    wire  [5 :0]  cp0_rtu_ex1_wb_preg,
  input    wire          cp0_rtu_ex1_wb_vld,
  input    wire          cp0_rtu_fence_idle,
  input    wire          cp0_rtu_icg_en,
  input    wire          cp0_rtu_in_lpmd,
  input    wire  [14:0]  cp0_rtu_int_vld,
  input    wire  [2 :0]  cp0_rtu_ecfg_vs,
  input    wire  [63:0]  cp0_rtu_trap_pc,
  input    wire          cp0_rtu_vstart_eq_0,
  input    wire          cp0_yy_clk_en,
  input    wire          cpurst_b,
  input    wire          dtu_rtu_async_halt_req,
  input    wire  [63:0]  dtu_rtu_dpc,
  input    wire          dtu_rtu_ebreak_action,
  input    wire          dtu_rtu_int_mask,
  input    wire  [63:0]  dtu_rtu_pending_tval,
  input    wire          dtu_rtu_resume_req,
  input    wire          dtu_rtu_step_en,
  input    wire          dtu_rtu_sync_flush,
  input    wire          dtu_rtu_sync_halt_req,
  input    wire          forever_cpuclk,
  input    wire          hpcp_rtu_cnt_en,
  input    wire          ifu_rtu_reset_halt_req,
  input    wire          ifu_rtu_warm_up,
  input    wire          iu_rtu_depd_lsu_chgflow_vld,
  input    wire  [63:0]  iu_rtu_depd_lsu_next_pc,
  input    wire  [63:0]  iu_rtu_div_data,
  input    wire  [5 :0]  iu_rtu_div_preg,
  input    wire          iu_rtu_div_wb_dp,
  input    wire          iu_rtu_div_wb_vld,
  input    wire          iu_rtu_ex1_alu_cmplt,
  input    wire          iu_rtu_ex1_alu_cmplt_dp,
  input    wire  [63:0]  iu_rtu_ex1_alu_data,
  input    wire          iu_rtu_ex1_alu_inst_len,
  input    wire          iu_rtu_ex1_alu_inst_split,
  input    wire  [5 :0]  iu_rtu_ex1_alu_preg,
  input    wire          iu_rtu_ex1_alu_wb_dp,
  input    wire          iu_rtu_ex1_alu_wb_vld,
  input    wire          iu_rtu_ex1_bju_cmplt,
  input    wire          iu_rtu_ex1_bju_cmplt_dp,
  input    wire  [63:0]  iu_rtu_ex1_bju_data,
  input    wire          iu_rtu_ex1_bju_inst_len,
  input    wire  [5 :0]  iu_rtu_ex1_bju_preg,
  input    wire          iu_rtu_ex1_bju_wb_dp,
  input    wire          iu_rtu_ex1_bju_wb_vld,
  input    wire          iu_rtu_ex1_branch_inst,
  input    wire  [63:0]  iu_rtu_ex1_cur_pc,
  input    wire          iu_rtu_ex1_div_cmplt,
  input    wire          iu_rtu_ex1_div_cmplt_dp,
  input    wire          iu_rtu_ex1_mul_cmplt,
  input    wire          iu_rtu_ex1_mul_cmplt_dp,
  input    wire  [63:0]  iu_rtu_ex1_next_pc,
  input    wire          iu_rtu_ex2_bju_ras_mispred,
  input    wire  [63:0]  iu_rtu_ex3_mul_data,
  input    wire  [5 :0]  iu_rtu_ex3_mul_preg,
  input    wire          iu_rtu_ex3_mul_wb_vld,
  input    wire          iu_xx_no_op,
  input    wire          lsu_rtu_async_expt_vld,
  input    wire          lsu_rtu_async_ld_inst,
  input    wire  [39:0]  lsu_rtu_async_tval,
  input    wire          lsu_rtu_ex1_buffer_vld,
  input    wire          lsu_rtu_ex1_cmplt,
  input    wire          lsu_rtu_ex1_cmplt_dp,
  input    wire          lsu_rtu_ex1_cmplt_for_pcgen,
  input    wire  [63:0]  lsu_rtu_ex1_data,
  input    wire  [5 :0]  lsu_rtu_ex1_dest_reg,
  input    wire  [39:0]  lsu_rtu_ex1_expt_tval,
  input    wire  [14:0]  lsu_rtu_ex1_expt_vec,
  input    wire          lsu_rtu_ex1_expt_vld,
  input    wire          lsu_rtu_ex1_fs_dirty,
  input    wire  [21:0]  lsu_rtu_ex1_halt_info,
  input    wire          lsu_rtu_ex1_inst_len,
  input    wire          lsu_rtu_ex1_inst_split,
  input    wire          lsu_rtu_ex1_tval2_vld,
  input    wire          lsu_rtu_ex1_vs_dirty,
  input    wire  [6 :0]  lsu_rtu_ex1_vstart,
  input    wire          lsu_rtu_ex1_vstart_vld,
  input    wire          lsu_rtu_ex1_wb_dp,
  input    wire          lsu_rtu_ex1_wb_vld,
  input    wire  [63:0]  lsu_rtu_ex2_data,
  input    wire          lsu_rtu_ex2_data_vld,
  input    wire  [5 :0]  lsu_rtu_ex2_dest_reg,
  input    wire  [39:0]  lsu_rtu_ex2_tval2,
  input    wire          lsu_rtu_no_op,
  input    wire  [63:0]  lsu_rtu_wb_data,
  input    wire  [5 :0]  lsu_rtu_wb_dest_reg,
  input    wire          lsu_rtu_wb_vld,
  input    wire          mmu_xx_mmu_en,
  input    wire          pad_yy_icg_scan_en,
  input    wire          vidu_rtu_no_op,
  input    wire  [7 :0]  vlsu_rtu_vl_updt_data,
  input    wire          vlsu_rtu_vl_updt_vld,
  input    wire          vpu_rtu_ex1_cmplt,
  input    wire          vpu_rtu_ex1_cmplt_dp,
  input    wire          vpu_rtu_ex1_inst_split,
  input    wire          vpu_rtu_ex1_fp_dirty,
  input    wire          vpu_rtu_ex1_vec_dirty,
  input    wire  [5 :0]  vpu_rtu_fflag,
  input    wire          vpu_rtu_fflag_vld,
  input    wire  [1 :0]  vpu_rtu_fflag_num,
  input    wire          vpu_rtu_split_vld,
  input    wire  [63:0]  vpu_rtu_gpr_wb_data,
  input    wire  [5 :0]  vpu_rtu_gpr_wb_index,
  input    wire          vpu_rtu_gpr_wb_req,
  input    wire          vpu_rtu_fcc_wb_req,
  input    wire  [2 :0]  vpu_rtu_fcc_wb_index,
  input    wire          vpu_rtu_fcc_wb_data,
  input    wire          vpu_rtu_no_op,
  input    wire          vpu_rtu_inst_expt_vld,
  output   wire  [63:0]  rtu_cp0_epc,
  output   wire          rtu_cp0_exit_debug,
  output   wire  [4 :0]  rtu_cp0_fflags,
  output   wire          rtu_cp0_fflags_updt,
  output   wire          rtu_cp0_split_vld,
  output   wire          rtu_cp0_fs_dirty_updt,
  output   wire          rtu_cp0_fs_dirty_updt_dp,
  output   wire  [63:0]  rtu_cp0_tval,
  output   wire  [7 :0]  rtu_cp0_vl,
  output   wire          rtu_cp0_vl_vld,
  output   wire          rtu_cp0_vs_dirty_updt,
  output   wire          rtu_cp0_vs_dirty_updt_dp,
  output   wire  [6 :0]  rtu_cp0_vstart,
  output   wire          rtu_cp0_vstart_vld,
  output   wire          rtu_cp0_vxsat,
  output   wire          rtu_cp0_vxsat_vld,
  output   wire          rtu_cpu_no_retire,
  output   wire  [14:0]  rtu_dtu_debug_info,
  output   wire  [63:0]  rtu_dtu_dpc,
  output   wire          rtu_dtu_halt_ack,
  output   wire          rtu_dtu_pending_ack,
  output   wire          rtu_dtu_retire_chgflw,
  output   wire          rtu_dtu_retire_debug_expt_vld,
  output   wire  [21:0]  rtu_dtu_retire_halt_info,
  output   wire          rtu_dtu_retire_ertn,
  output   wire          rtu_dtu_retire_mret,
  output   wire  [63:0]  rtu_dtu_retire_next_pc,
  output   wire          rtu_dtu_retire_sret,
  output   wire          rtu_dtu_retire_vld,
  output   wire  [63:0]  rtu_dtu_tval,
  output   wire          rtu_hpcp_int_vld,
  output   wire          rtu_hpcp_retire_inst_vld,
  output   wire  [63:0]  rtu_hpcp_retire_pc,
  output   wire          rtu_idu_commit,
  output   wire          rtu_idu_commit_for_bju,
  output   wire          rtu_idu_flush_fe,
  output   wire          rtu_idu_flush_stall,
  output   wire          rtu_idu_flush_wbt,
  output   wire  [63:0]  rtu_idu_fwd0_data,
  output   wire  [5 :0]  rtu_idu_fwd0_reg,
  output   wire          rtu_idu_fwd0_vld,
  output   wire  [63:0]  rtu_idu_fwd1_data,
  output   wire  [5 :0]  rtu_idu_fwd1_reg,
  output   wire          rtu_idu_fwd1_vld,
  output   wire  [63:0]  rtu_idu_fwd2_data,
  output   wire  [5 :0]  rtu_idu_fwd2_reg,
  output   wire          rtu_idu_fwd2_vld,
  output   wire          rtu_idu_pipeline_empty,
  output   wire  [63:0]  rtu_idu_wb0_data,
  output   wire  [5 :0]  rtu_idu_wb0_reg,
  output   wire          rtu_idu_wb0_vld,
  output   wire  [63:0]  rtu_idu_wb1_data,
  output   wire  [5 :0]  rtu_idu_wb1_reg,
  output   wire          rtu_idu_wb1_vld,
  output   wire          rtu_idu_wbc_data,
  output   wire  [2 :0]  rtu_idu_wbc_reg,
  output   wire          rtu_idu_wbc_vld,
  output   wire          rtu_idu_wbe_vld,
  output   wire  [1 :0]  rtu_idu_wbe_num,
  output   wire  [63:0]  rtu_ifu_chgflw_pc,
  output   wire          rtu_ifu_chgflw_vld,
  output   wire          rtu_ifu_dbg_mask,
  output   wire          rtu_ifu_flush_fe,
  output   wire          rtu_iu_div_wb_grant,
  output   wire          rtu_iu_div_wb_grant_for_full,
  output   wire          rtu_iu_ex1_cmplt,
  output   wire          rtu_iu_ex1_cmplt_dp,
  output   wire          rtu_iu_ex1_inst_len,
  output   wire          rtu_iu_ex1_inst_split,
  output   wire  [63:0]  rtu_iu_ex2_cur_pc,
  output   wire  [63:0]  rtu_iu_ex2_next_pc,
  output   wire          rtu_iu_mul_wb_grant,
  output   wire          rtu_iu_mul_wb_grant_for_full,
  output   wire          rtu_lsu_async_expt_ack,
  output   wire          rtu_lsu_expt_ack,
  output   wire          rtu_lsu_expt_exit,
  output   wire  [26:0]  rtu_mmu_bad_vpn,
  output   wire          rtu_mmu_expt_vld,
  output   wire          rtu_pad_halted,
  output   wire          rtu_pad_retire,
  output   wire  [63:0]  rtu_pad_retire_pc,
  output   wire          rtu_vidu_flush_wbt,
  output   wire          rtu_vpu_gpr_wb_grnt,
  output   wire          rtu_yy_xx_async_flush,
  output   wire          rtu_yy_xx_dbgon,
  output   wire          rtu_yy_xx_expt_int,
  output   wire  [14:0]  rtu_yy_xx_expt_vec,
  output   wire          rtu_yy_xx_expt_vld,
  output   wire          rtu_yy_xx_flush,
  output   wire          rtu_yy_xx_flush_fe
); 



// &Regs; @26
// &Wires; @27
wire            async_select_next_pc;            
wire            ctrl_dp_ex1_cmplt_dp;            
wire            ctrl_retire_ex2_retire_vld;      
wire            ctrl_top_dbg_info;               
wire            dp_ctrl_ex1_cmplt_dp;            
wire            dp_int_ex2_inst_split;           
wire            dp_misc_clk;                     
wire    [63:0]  dp_retire_ex2_cur_pc;            
wire            dp_retire_ex2_fs_dirty;          
wire    [21:0]  dp_retire_ex2_halt_info;         
wire            dp_retire_ex2_inst_branch;       
wire            dp_retire_ex2_inst_chgflw;       
wire            dp_retire_ex2_inst_dret;         
wire            dp_retire_ex2_inst_ebreak;       
wire            dp_retire_ex2_inst_expt;         
wire            dp_retire_ex2_inst_flush;        
wire            dp_retire_ex2_inst_mret;         
wire            dp_retire_ex2_inst_split;        
wire            dp_retire_ex2_inst_sret;         
wire            dp_retire_ex2_inst_vstart;       
wire    [63:0]  dp_retire_ex2_next_pc;           
wire    [63:0]  dp_retire_ex2_tval;              
wire    [14:0]  dp_retire_ex2_vec;               
wire            dp_retire_ex2_vs_dirty;          
wire    [6 :0]  dp_retire_ex2_vstart;            
wire    [2 :0]  dp_top_dbg_info;                 
wire    [14:0]  int_retire_int_vec;              
wire            int_retire_int_vld;              
wire    [63:0]  rbus_wb_rbus_wb_data;            
wire            rbus_wb_rbus_wb_dp;              
wire    [5 :0]  rbus_wb_rbus_wb_preg;            
wire            rbus_wb_rbus_wb_vld;             
wire            retire_ctrl_commit_clear;        
wire            retire_ctrl_commit_clear_for_bju; 
wire            retire_rbus_fs_dirty;            
wire            retire_rbus_vs_dirty;            
wire    [10:0]  retire_top_dbg_info;             
wire            wb_retire_wb_no_op;              


// &Instance("aq_rtu_ctrl"); @29
aq_rtu_ctrl  x_aq_rtu_ctrl (
  .async_select_next_pc             (async_select_next_pc            ),
  .cp0_rtu_ex1_cmplt                (cp0_rtu_ex1_cmplt               ),
  .cp0_rtu_icg_en                   (cp0_rtu_icg_en                  ),
  .cp0_yy_clk_en                    (cp0_yy_clk_en                   ),
  .cpurst_b                         (cpurst_b                        ),
  .ctrl_dp_ex1_cmplt_dp             (ctrl_dp_ex1_cmplt_dp            ),
  .ctrl_retire_ex2_retire_vld       (ctrl_retire_ex2_retire_vld      ),
  .ctrl_top_dbg_info                (ctrl_top_dbg_info               ),
  .dp_ctrl_ex1_cmplt_dp             (dp_ctrl_ex1_cmplt_dp            ),
  .dp_misc_clk                      (dp_misc_clk                     ),
  .forever_cpuclk                   (forever_cpuclk                  ),
  .ifu_rtu_warm_up                  (ifu_rtu_warm_up                 ),
  .iu_rtu_ex1_alu_cmplt             (iu_rtu_ex1_alu_cmplt            ),
  .iu_rtu_ex1_bju_cmplt             (iu_rtu_ex1_bju_cmplt            ),
  .iu_rtu_ex1_div_cmplt             (iu_rtu_ex1_div_cmplt            ),
  .iu_rtu_ex1_mul_cmplt             (iu_rtu_ex1_mul_cmplt            ),
  .lsu_rtu_ex1_cmplt                (lsu_rtu_ex1_cmplt               ),
  .lsu_rtu_ex1_cmplt_for_pcgen      (lsu_rtu_ex1_cmplt_for_pcgen     ),
  .pad_yy_icg_scan_en               (pad_yy_icg_scan_en              ),
  .retire_ctrl_commit_clear         (retire_ctrl_commit_clear        ),
  .retire_ctrl_commit_clear_for_bju (retire_ctrl_commit_clear_for_bju),
  .rtu_idu_commit                   (rtu_idu_commit                  ),
  .rtu_idu_commit_for_bju           (rtu_idu_commit_for_bju          ),
  .rtu_iu_ex1_cmplt                 (rtu_iu_ex1_cmplt                ),
  .rtu_iu_ex1_cmplt_dp              (rtu_iu_ex1_cmplt_dp             ),
  .vpu_rtu_ex1_cmplt                (vpu_rtu_ex1_cmplt               )
);


// &Instance("aq_rtu_dp"); @31
aq_rtu_dp  x_aq_rtu_dp (
  .cp0_rtu_ex1_chgflw          (cp0_rtu_ex1_chgflw         ),
  .cp0_rtu_ex1_chgflw_pc       (cp0_rtu_ex1_chgflw_pc      ),
  .cp0_rtu_ex1_cmplt_dp        (cp0_rtu_ex1_cmplt_dp       ),
  .cp0_rtu_ex1_expt_tval       (cp0_rtu_ex1_expt_tval      ),
  .cp0_rtu_ex1_expt_vec        (cp0_rtu_ex1_expt_vec       ),
  .cp0_rtu_ex1_expt_vld        (cp0_rtu_ex1_expt_vld       ),
  .cp0_rtu_ex1_flush           (cp0_rtu_ex1_flush          ),
  .cp0_rtu_ex1_halt_info       (cp0_rtu_ex1_halt_info      ),
  .cp0_rtu_ex1_inst_dret       (cp0_rtu_ex1_inst_dret      ),
  .cp0_rtu_ex1_inst_ebreak     (cp0_rtu_ex1_inst_ebreak    ),
  .cp0_rtu_ex1_inst_len        (cp0_rtu_ex1_inst_len       ),
  .cp0_rtu_ex1_inst_ertn       (cp0_rtu_ex1_inst_ertn      ),
  .cp0_rtu_ex1_inst_mret       (cp0_rtu_ex1_inst_mret      ),
  .cp0_rtu_ex1_inst_split      (cp0_rtu_ex1_inst_split     ),
  .cp0_rtu_ex1_inst_sret       (cp0_rtu_ex1_inst_sret      ),
  .cp0_rtu_icg_en              (cp0_rtu_icg_en             ),
  .cp0_yy_clk_en               (cp0_yy_clk_en              ),
  .ctrl_dp_ex1_cmplt_dp        (ctrl_dp_ex1_cmplt_dp       ),
  .dp_ctrl_ex1_cmplt_dp        (dp_ctrl_ex1_cmplt_dp       ),
  .dp_int_ex2_inst_split       (dp_int_ex2_inst_split      ),
  .dp_misc_clk                 (dp_misc_clk                ),
  .dp_retire_ex2_cur_pc        (dp_retire_ex2_cur_pc       ),
  .dp_retire_ex2_fs_dirty      (dp_retire_ex2_fs_dirty     ),
  .dp_retire_ex2_halt_info     (dp_retire_ex2_halt_info    ),
  .dp_retire_ex2_inst_branch   (dp_retire_ex2_inst_branch  ),
  .dp_retire_ex2_inst_chgflw   (dp_retire_ex2_inst_chgflw  ),
  .dp_retire_ex2_inst_dret     (dp_retire_ex2_inst_dret    ),
  .dp_retire_ex2_inst_ebreak   (dp_retire_ex2_inst_ebreak  ),
  .dp_retire_ex2_inst_expt     (dp_retire_ex2_inst_expt    ),
  .dp_retire_ex2_inst_flush    (dp_retire_ex2_inst_flush   ),
  .dp_retire_ex2_inst_ertn     (dp_retire_ex2_inst_ertn    ),
  .dp_retire_ex2_inst_mret     (dp_retire_ex2_inst_mret    ),
  .dp_retire_ex2_inst_split    (dp_retire_ex2_inst_split   ),
  .dp_retire_ex2_inst_sret     (dp_retire_ex2_inst_sret    ),
  .dp_retire_ex2_inst_vstart   (dp_retire_ex2_inst_vstart  ),
  .dp_retire_ex2_next_pc       (dp_retire_ex2_next_pc      ),
  .dp_retire_ex2_tval          (dp_retire_ex2_tval         ),
  .dp_retire_ex2_vec           (dp_retire_ex2_vec          ),
  .dp_retire_ex2_vs_dirty      (dp_retire_ex2_vs_dirty     ),
  .dp_retire_ex2_vstart        (dp_retire_ex2_vstart       ),
  .dp_top_dbg_info             (dp_top_dbg_info            ),
  .forever_cpuclk              (forever_cpuclk             ),
  .ifu_rtu_warm_up             (ifu_rtu_warm_up            ),
  .iu_rtu_depd_lsu_chgflow_vld (iu_rtu_depd_lsu_chgflow_vld),
  .iu_rtu_depd_lsu_next_pc     (iu_rtu_depd_lsu_next_pc    ),
  .iu_rtu_ex1_alu_cmplt_dp     (iu_rtu_ex1_alu_cmplt_dp    ),
  .iu_rtu_ex1_alu_inst_len     (iu_rtu_ex1_alu_inst_len    ),
  .iu_rtu_ex1_alu_inst_split   (iu_rtu_ex1_alu_inst_split  ),
  .iu_rtu_ex1_bju_cmplt_dp     (iu_rtu_ex1_bju_cmplt_dp    ),
  .iu_rtu_ex1_bju_inst_len     (iu_rtu_ex1_bju_inst_len    ),
  .iu_rtu_ex1_branch_inst      (iu_rtu_ex1_branch_inst     ),
  .iu_rtu_ex1_cur_pc           (iu_rtu_ex1_cur_pc          ),
  .iu_rtu_ex1_div_cmplt_dp     (iu_rtu_ex1_div_cmplt_dp    ),
  .iu_rtu_ex1_mul_cmplt_dp     (iu_rtu_ex1_mul_cmplt_dp    ),
  .iu_rtu_ex1_next_pc          (iu_rtu_ex1_next_pc         ),
  .lsu_rtu_ex1_cmplt_dp        (lsu_rtu_ex1_cmplt_dp       ),
  .lsu_rtu_ex1_expt_tval       (lsu_rtu_ex1_expt_tval      ),
  .lsu_rtu_ex1_expt_vec        (lsu_rtu_ex1_expt_vec       ),
  .lsu_rtu_ex1_expt_vld        (lsu_rtu_ex1_expt_vld       ),
  .lsu_rtu_ex1_fs_dirty        (lsu_rtu_ex1_fs_dirty       ),
  .lsu_rtu_ex1_halt_info       (lsu_rtu_ex1_halt_info      ),
  .lsu_rtu_ex1_inst_len        (lsu_rtu_ex1_inst_len       ),
  .lsu_rtu_ex1_inst_split      (lsu_rtu_ex1_inst_split     ),
  .lsu_rtu_ex1_tval2_vld       (lsu_rtu_ex1_tval2_vld      ),
  .lsu_rtu_ex1_vs_dirty        (lsu_rtu_ex1_vs_dirty       ),
  .lsu_rtu_ex1_vstart          (lsu_rtu_ex1_vstart         ),
  .lsu_rtu_ex1_vstart_vld      (lsu_rtu_ex1_vstart_vld     ),
  .lsu_rtu_ex2_tval2           (lsu_rtu_ex2_tval2          ),
  .pad_yy_icg_scan_en          (pad_yy_icg_scan_en         ),
  .rtu_iu_ex1_inst_len         (rtu_iu_ex1_inst_len        ),
  .rtu_iu_ex1_inst_split       (rtu_iu_ex1_inst_split      ),
  .rtu_iu_ex2_cur_pc           (rtu_iu_ex2_cur_pc          ),
  .rtu_iu_ex2_next_pc          (rtu_iu_ex2_next_pc         ),
  .vpu_rtu_ex1_cmplt_dp        (vpu_rtu_ex1_cmplt_dp       ),
  .vpu_rtu_ex1_inst_split      (vpu_rtu_ex1_inst_split     ),
  .vpu_rtu_inst_expt_vld       (vpu_rtu_inst_expt_vld      )
);


// &Instance("aq_rtu_rbus"); @33
aq_rtu_rbus  x_aq_rtu_rbus (
  .forever_cpuclk               (forever_cpuclk              ),
  .cpurst_b                     (cpurst_b                    ),
  .cp0_rtu_ex1_cmplt            (cp0_rtu_ex1_cmplt           ),
  .cp0_rtu_ex1_cmplt_dp         (cp0_rtu_ex1_cmplt_dp        ),
  .cp0_rtu_ex1_vs_dirty         (cp0_rtu_ex1_vs_dirty        ),
  .cp0_rtu_ex1_vs_dirty_dp      (cp0_rtu_ex1_vs_dirty_dp     ),
  .cp0_rtu_ex1_wb_data          (cp0_rtu_ex1_wb_data         ),
  .cp0_rtu_ex1_wb_dp            (cp0_rtu_ex1_wb_dp           ),
  .cp0_rtu_ex1_wb_preg          (cp0_rtu_ex1_wb_preg         ),
  .cp0_rtu_ex1_wb_vld           (cp0_rtu_ex1_wb_vld          ),
  .iu_rtu_div_data              (iu_rtu_div_data             ),
  .iu_rtu_div_preg              (iu_rtu_div_preg             ),
  .iu_rtu_div_wb_dp             (iu_rtu_div_wb_dp            ),
  .iu_rtu_div_wb_vld            (iu_rtu_div_wb_vld           ),
  .iu_rtu_ex1_alu_data          (iu_rtu_ex1_alu_data         ),
  .iu_rtu_ex1_alu_preg          (iu_rtu_ex1_alu_preg         ),
  .iu_rtu_ex1_alu_wb_dp         (iu_rtu_ex1_alu_wb_dp        ),
  .iu_rtu_ex1_alu_wb_vld        (iu_rtu_ex1_alu_wb_vld       ),
  .iu_rtu_ex1_bju_data          (iu_rtu_ex1_bju_data         ),
  .iu_rtu_ex1_bju_preg          (iu_rtu_ex1_bju_preg         ),
  .iu_rtu_ex1_bju_wb_dp         (iu_rtu_ex1_bju_wb_dp        ),
  .iu_rtu_ex1_bju_wb_vld        (iu_rtu_ex1_bju_wb_vld       ),
  .iu_rtu_ex3_mul_data          (iu_rtu_ex3_mul_data         ),
  .iu_rtu_ex3_mul_preg          (iu_rtu_ex3_mul_preg         ),
  .iu_rtu_ex3_mul_wb_vld        (iu_rtu_ex3_mul_wb_vld       ),
  .lsu_rtu_ex1_data             (lsu_rtu_ex1_data            ),
  .lsu_rtu_ex1_dest_reg         (lsu_rtu_ex1_dest_reg        ),
  .lsu_rtu_ex1_wb_dp            (lsu_rtu_ex1_wb_dp           ),
  .lsu_rtu_ex1_wb_vld           (lsu_rtu_ex1_wb_vld          ),
  .lsu_rtu_ex2_data             (lsu_rtu_ex2_data            ),
  .lsu_rtu_ex2_data_vld         (lsu_rtu_ex2_data_vld        ),
  .lsu_rtu_ex2_dest_reg         (lsu_rtu_ex2_dest_reg        ),
  .rtu_pad_retire               (rtu_pad_retire              ),
  .rtu_pad_retire_pc            (rtu_pad_retire_pc           ),
  .rbus_wb_rbus_wb_data         (rbus_wb_rbus_wb_data        ),
  .rbus_wb_rbus_wb_dp           (rbus_wb_rbus_wb_dp          ),
  .rbus_wb_rbus_wb_preg         (rbus_wb_rbus_wb_preg        ),
  .rbus_wb_rbus_wb_vld          (rbus_wb_rbus_wb_vld         ),
  .retire_rbus_fs_dirty         (retire_rbus_fs_dirty        ),
  .retire_rbus_vs_dirty         (retire_rbus_vs_dirty        ),
  .rtu_cp0_fs_dirty_updt        (rtu_cp0_fs_dirty_updt       ),
  .rtu_cp0_fs_dirty_updt_dp     (rtu_cp0_fs_dirty_updt_dp    ),
  .rtu_cp0_vl                   (rtu_cp0_vl                  ),
  .rtu_cp0_vl_vld               (rtu_cp0_vl_vld              ),
  .rtu_cp0_vs_dirty_updt        (rtu_cp0_vs_dirty_updt       ),
  .rtu_cp0_vs_dirty_updt_dp     (rtu_cp0_vs_dirty_updt_dp    ),
  .rtu_idu_fwd0_data            (rtu_idu_fwd0_data           ),
  .rtu_idu_fwd0_reg             (rtu_idu_fwd0_reg            ),
  .rtu_idu_fwd0_vld             (rtu_idu_fwd0_vld            ),
  .rtu_idu_fwd1_data            (rtu_idu_fwd1_data           ),
  .rtu_idu_fwd1_reg             (rtu_idu_fwd1_reg            ),
  .rtu_idu_fwd1_vld             (rtu_idu_fwd1_vld            ),
  .rtu_idu_fwd2_data            (rtu_idu_fwd2_data           ),
  .rtu_idu_fwd2_reg             (rtu_idu_fwd2_reg            ),
  .rtu_idu_fwd2_vld             (rtu_idu_fwd2_vld            ),
  .rtu_iu_div_wb_grant          (rtu_iu_div_wb_grant         ),
  .rtu_iu_div_wb_grant_for_full (rtu_iu_div_wb_grant_for_full),
  .rtu_iu_mul_wb_grant          (rtu_iu_mul_wb_grant         ),
  .rtu_iu_mul_wb_grant_for_full (rtu_iu_mul_wb_grant_for_full),
  .vlsu_rtu_vl_updt_data        (vlsu_rtu_vl_updt_data       ),
  .vlsu_rtu_vl_updt_vld         (vlsu_rtu_vl_updt_vld        ),
  .vpu_rtu_ex1_cmplt            (vpu_rtu_ex1_cmplt           ),
  .vpu_rtu_ex1_cmplt_dp         (vpu_rtu_ex1_cmplt_dp        ),
  .vpu_rtu_ex1_fp_dirty         (vpu_rtu_ex1_fp_dirty        ),
  .vpu_rtu_ex1_vec_dirty        (vpu_rtu_ex1_vec_dirty       )
);


// &Instance("aq_rtu_retire"); @35
aq_rtu_retire  x_aq_rtu_retire (
  .async_select_next_pc             (async_select_next_pc            ),
  .cp0_rtu_fence_idle               (cp0_rtu_fence_idle              ),
  .cp0_rtu_icg_en                   (cp0_rtu_icg_en                  ),
  .cp0_rtu_in_lpmd                  (cp0_rtu_in_lpmd                 ),
  .cp0_rtu_trap_pc                  (cp0_rtu_trap_pc                 ),
  .cp0_rtu_vstart_eq_0              (cp0_rtu_vstart_eq_0             ),
  .cp0_yy_clk_en                    (cp0_yy_clk_en                   ),
  .cpurst_b                         (cpurst_b                        ),
  .ctrl_retire_ex2_retire_vld       (ctrl_retire_ex2_retire_vld      ),
  .dp_retire_ex2_cur_pc             (dp_retire_ex2_cur_pc            ),
  .dp_retire_ex2_fs_dirty           (dp_retire_ex2_fs_dirty          ),
  .dp_retire_ex2_halt_info          (dp_retire_ex2_halt_info         ),
  .dp_retire_ex2_inst_branch        (dp_retire_ex2_inst_branch       ),
  .dp_retire_ex2_inst_chgflw        (dp_retire_ex2_inst_chgflw       ),
  .dp_retire_ex2_inst_dret          (dp_retire_ex2_inst_dret         ),
  .dp_retire_ex2_inst_ebreak        (dp_retire_ex2_inst_ebreak       ),
  .dp_retire_ex2_inst_expt          (dp_retire_ex2_inst_expt         ),
  .dp_retire_ex2_inst_flush         (dp_retire_ex2_inst_flush        ),
  .dp_retire_ex2_inst_ertn          (dp_retire_ex2_inst_ertn         ),
  .dp_retire_ex2_inst_mret          (dp_retire_ex2_inst_mret         ),
  .dp_retire_ex2_inst_split         (dp_retire_ex2_inst_split        ),
  .dp_retire_ex2_inst_sret          (dp_retire_ex2_inst_sret         ),
  .dp_retire_ex2_inst_vstart        (dp_retire_ex2_inst_vstart       ),
  .dp_retire_ex2_next_pc            (dp_retire_ex2_next_pc           ),
  .dp_retire_ex2_tval               (dp_retire_ex2_tval              ),
  .dp_retire_ex2_vec                (dp_retire_ex2_vec               ),
  .dp_retire_ex2_vs_dirty           (dp_retire_ex2_vs_dirty          ),
  .dp_retire_ex2_vstart             (dp_retire_ex2_vstart            ),
  .dtu_rtu_async_halt_req           (dtu_rtu_async_halt_req          ),
  .dtu_rtu_dpc                      (dtu_rtu_dpc                     ),
  .dtu_rtu_ebreak_action            (dtu_rtu_ebreak_action           ),
  .dtu_rtu_pending_tval             (dtu_rtu_pending_tval            ),
  .dtu_rtu_resume_req               (dtu_rtu_resume_req              ),
  .dtu_rtu_step_en                  (dtu_rtu_step_en                 ),
  .dtu_rtu_sync_flush               (dtu_rtu_sync_flush              ),
  .dtu_rtu_sync_halt_req            (dtu_rtu_sync_halt_req           ),
  .forever_cpuclk                   (forever_cpuclk                  ),
  .hpcp_rtu_cnt_en                  (hpcp_rtu_cnt_en                 ),
  .ifu_rtu_reset_halt_req           (ifu_rtu_reset_halt_req          ),
  .ifu_rtu_warm_up                  (ifu_rtu_warm_up                 ),
  .int_retire_int_vec               (int_retire_int_vec              ),
  .int_retire_int_vld               (int_retire_int_vld              ),
  .iu_rtu_depd_lsu_chgflow_vld      (iu_rtu_depd_lsu_chgflow_vld     ),
  .iu_rtu_ex2_bju_ras_mispred       (iu_rtu_ex2_bju_ras_mispred      ),
  .iu_xx_no_op                      (iu_xx_no_op                     ),
  .lsu_rtu_async_expt_vld           (lsu_rtu_async_expt_vld          ),
  .lsu_rtu_async_ld_inst            (lsu_rtu_async_ld_inst           ),
  .lsu_rtu_async_tval               (lsu_rtu_async_tval              ),
  .lsu_rtu_ex1_buffer_vld           (lsu_rtu_ex1_buffer_vld          ),
  .lsu_rtu_no_op                    (lsu_rtu_no_op                   ),
  .mmu_xx_mmu_en                    (mmu_xx_mmu_en                   ),
  .pad_yy_icg_scan_en               (pad_yy_icg_scan_en              ),
  .retire_ctrl_commit_clear         (retire_ctrl_commit_clear        ),
  .retire_ctrl_commit_clear_for_bju (retire_ctrl_commit_clear_for_bju),
  .retire_rbus_fs_dirty             (retire_rbus_fs_dirty            ),
  .retire_rbus_vs_dirty             (retire_rbus_vs_dirty            ),
  .retire_top_dbg_info              (retire_top_dbg_info             ),
  .rtu_cp0_epc                      (rtu_cp0_epc                     ),
  .rtu_cp0_exit_debug               (rtu_cp0_exit_debug              ),
  .rtu_cp0_tval                     (rtu_cp0_tval                    ),
  .rtu_cp0_vstart                   (rtu_cp0_vstart                  ),
  .rtu_cp0_vstart_vld               (rtu_cp0_vstart_vld              ),
  .rtu_cpu_no_retire                (rtu_cpu_no_retire               ),
  .rtu_dtu_dpc                      (rtu_dtu_dpc                     ),
  .rtu_dtu_halt_ack                 (rtu_dtu_halt_ack                ),
  .rtu_dtu_pending_ack              (rtu_dtu_pending_ack             ),
  .rtu_dtu_retire_chgflw            (rtu_dtu_retire_chgflw           ),
  .rtu_dtu_retire_debug_expt_vld    (rtu_dtu_retire_debug_expt_vld   ),
  .rtu_dtu_retire_halt_info         (rtu_dtu_retire_halt_info        ),
  .rtu_dtu_retire_ertn              (rtu_dtu_retire_ertn             ),
  .rtu_dtu_retire_mret              (rtu_dtu_retire_mret             ),
  .rtu_dtu_retire_next_pc           (rtu_dtu_retire_next_pc          ),
  .rtu_dtu_retire_sret              (rtu_dtu_retire_sret             ),
  .rtu_dtu_retire_vld               (rtu_dtu_retire_vld              ),
  .rtu_dtu_tval                     (rtu_dtu_tval                    ),
  .rtu_hpcp_int_vld                 (rtu_hpcp_int_vld                ),
  .rtu_hpcp_retire_inst_vld         (rtu_hpcp_retire_inst_vld        ),
  .rtu_hpcp_retire_pc               (rtu_hpcp_retire_pc              ),
  .rtu_idu_flush_fe                 (rtu_idu_flush_fe                ),
  .rtu_idu_flush_stall              (rtu_idu_flush_stall             ),
  .rtu_idu_flush_wbt                (rtu_idu_flush_wbt               ),
  .rtu_idu_pipeline_empty           (rtu_idu_pipeline_empty          ),
  .rtu_ifu_chgflw_pc                (rtu_ifu_chgflw_pc               ),
  .rtu_ifu_chgflw_vld               (rtu_ifu_chgflw_vld              ),
  .rtu_ifu_dbg_mask                 (rtu_ifu_dbg_mask                ),
  .rtu_ifu_flush_fe                 (rtu_ifu_flush_fe                ),
  .rtu_lsu_async_expt_ack           (rtu_lsu_async_expt_ack          ),
  .rtu_lsu_expt_ack                 (rtu_lsu_expt_ack                ),
  .rtu_lsu_expt_exit                (rtu_lsu_expt_exit               ),
  .rtu_mmu_bad_vpn                  (rtu_mmu_bad_vpn                 ),
  .rtu_mmu_expt_vld                 (rtu_mmu_expt_vld                ),
  .rtu_pad_halted                   (rtu_pad_halted                  ),
  .rtu_pad_retire                   (rtu_pad_retire                  ),
  .rtu_pad_retire_pc                (rtu_pad_retire_pc               ),
  .rtu_vidu_flush_wbt               (rtu_vidu_flush_wbt              ),
  .rtu_yy_xx_async_flush            (rtu_yy_xx_async_flush           ),
  .rtu_yy_xx_dbgon                  (rtu_yy_xx_dbgon                 ),
  .rtu_yy_xx_expt_int               (rtu_yy_xx_expt_int              ),
  .rtu_yy_xx_expt_vec               (rtu_yy_xx_expt_vec              ),
  .rtu_yy_xx_expt_vld               (rtu_yy_xx_expt_vld              ),
  .rtu_yy_xx_flush                  (rtu_yy_xx_flush                 ),
  .rtu_yy_xx_flush_fe               (rtu_yy_xx_flush_fe              ),
  .vidu_rtu_no_op                   (vidu_rtu_no_op                  ),
  .vpu_rtu_no_op                    (vpu_rtu_no_op                   ),
  .wb_retire_wb_no_op               (wb_retire_wb_no_op              )
);


// &Instance("aq_rtu_wb"); @37
aq_rtu_wb  x_aq_rtu_wb (
  .cp0_rtu_icg_en       (cp0_rtu_icg_en      ),
  .cp0_yy_clk_en        (cp0_yy_clk_en       ),
  .cpurst_b             (cpurst_b            ),
  .forever_cpuclk       (forever_cpuclk      ),
  .ifu_rtu_warm_up      (ifu_rtu_warm_up     ),
  .lsu_rtu_wb_data      (lsu_rtu_wb_data     ),
  .lsu_rtu_wb_dest_reg  (lsu_rtu_wb_dest_reg ),
  .lsu_rtu_wb_vld       (lsu_rtu_wb_vld      ),
  .pad_yy_icg_scan_en   (pad_yy_icg_scan_en  ),
  .rbus_wb_rbus_wb_data (rbus_wb_rbus_wb_data),
  .rbus_wb_rbus_wb_dp   (rbus_wb_rbus_wb_dp  ),
  .rbus_wb_rbus_wb_preg (rbus_wb_rbus_wb_preg),
  .rbus_wb_rbus_wb_vld  (rbus_wb_rbus_wb_vld ),
  .rtu_cp0_fflags       (rtu_cp0_fflags      ),
  .rtu_cp0_fflags_updt  (rtu_cp0_fflags_updt ),
  .rtu_cp0_split_vld    (rtu_cp0_split_vld   ),
  .rtu_cp0_vxsat        (rtu_cp0_vxsat       ),
  .rtu_cp0_vxsat_vld    (rtu_cp0_vxsat_vld   ),
  .rtu_idu_wb0_data     (rtu_idu_wb0_data    ),
  .rtu_idu_wb0_reg      (rtu_idu_wb0_reg     ),
  .rtu_idu_wb0_vld      (rtu_idu_wb0_vld     ),
  .rtu_idu_wb1_data     (rtu_idu_wb1_data    ),
  .rtu_idu_wb1_reg      (rtu_idu_wb1_reg     ),
  .rtu_idu_wb1_vld      (rtu_idu_wb1_vld     ),
  .rtu_idu_wbc_data     (rtu_idu_wbc_data    ),
  .rtu_idu_wbc_reg      (rtu_idu_wbc_reg     ),
  .rtu_idu_wbc_vld      (rtu_idu_wbc_vld     ),
  .rtu_idu_wbe_vld      (rtu_idu_wbe_vld     ),
  .rtu_idu_wbe_num      (rtu_idu_wbe_num     ),
  .rtu_vpu_gpr_wb_grnt  (rtu_vpu_gpr_wb_grnt ),
  .vpu_rtu_fflag        (vpu_rtu_fflag       ),
  .vpu_rtu_fflag_vld    (vpu_rtu_fflag_vld   ),
  .vpu_rtu_fflag_num    (vpu_rtu_fflag_num   ),
  .vpu_rtu_split_vld    (vpu_rtu_split_vld   ),
  .vpu_rtu_gpr_wb_data  (vpu_rtu_gpr_wb_data ),
  .vpu_rtu_gpr_wb_index (vpu_rtu_gpr_wb_index),
  .vpu_rtu_gpr_wb_req   (vpu_rtu_gpr_wb_req  ),
  .vpu_rtu_fcc_wb_data  (vpu_rtu_fcc_wb_data ),
  .vpu_rtu_fcc_wb_index (vpu_rtu_fcc_wb_index),
  .vpu_rtu_fcc_wb_req   (vpu_rtu_fcc_wb_req  ),
  .wb_retire_wb_no_op   (wb_retire_wb_no_op  )
);


// &Instance("aq_rtu_int"); @39
aq_rtu_int  x_aq_rtu_int (
  .cp0_rtu_int_vld       (cp0_rtu_int_vld      ),
  .cp0_rtu_ecfg_vs       (cp0_rtu_ecfg_vs      ),
  .dp_int_ex2_inst_split (dp_int_ex2_inst_split),
  .dtu_rtu_int_mask      (dtu_rtu_int_mask     ),
  .int_retire_int_vec    (int_retire_int_vec   ),
  .int_retire_int_vld    (int_retire_int_vld   )
);


// &Force("output", "rtu_yy_xx_dbgon"); @41

assign rtu_dtu_debug_info[14:0] = {retire_top_dbg_info[10:0],
                                   ctrl_top_dbg_info,
                                   dp_top_dbg_info[2:0]};


// &ModuleEnd; @124
endmodule



