/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/
module ct_vfalu_top_pipe7 (
  // &Ports, @23
  input    wire          cp0_vfpu_icg_en,
  input    wire          cp0_yy_clk_en,
  input    wire          cpurst_b,
  input    wire  [19:0]  dp_vfalu_ex1_pipex_func,
  input    wire  [2 :0]  dp_vfalu_ex1_pipex_imm0,
  input    wire  [63:0]  dp_vfalu_ex1_pipex_mtvr_src0,
  input    wire  [2 :0]  dp_vfalu_ex1_pipex_sel,
  input    wire  [63:0]  dp_vfalu_ex1_pipex_srcf0,
  input    wire  [63:0]  dp_vfalu_ex1_pipex_srcf1,
  input    wire  [63:0]  dp_vfalu_ex1_pipex_srcf2,
  input    wire          forever_cpuclk,
  input    wire          pad_yy_icg_scan_en,
  input    wire          vfpu_yy_xx_dqnan,
  input    wire  [2 :0]  vfpu_yy_xx_rm,
  output   wire  [63:0]  pipex_dp_ex1_vfalu_mfvr_data,
  output   wire  [4 :0]  pipex_dp_ex3_vfalu_ereg_data,
  output   wire  [63:0]  pipex_dp_ex3_vfalu_freg_data
); 



// &Regs; @24
// &Wires; @25
wire            fadd_ereg_ex3_forward_r_vld; 
wire    [4 :0]  fadd_ereg_ex3_result;        
wire            fadd_forward_r_vld;          
wire    [63:0]  fadd_forward_result;         
wire    [63:0]  fadd_mfvr_cmp_result;        
wire            fcnvt_ereg_forward_r_vld;    
wire    [4 :0]  fcnvt_ereg_forward_result;   
wire            fcnvt_forward_r_vld;         
wire    [63:0]  fcnvt_forward_result;        
wire            fspu_forward_r_vld;          
wire    [63:0]  fspu_forward_result;         
wire    [63:0]  fspu_mfvr_data;              


// &Instance("ct_fcnvt_top"); @27
ct_fcnvt_top  x_ct_fcnvt_top (
  .cp0_vfpu_icg_en           (cp0_vfpu_icg_en          ),
  .cp0_yy_clk_en             (cp0_yy_clk_en            ),
  .cpurst_b                  (cpurst_b                 ),
  .dp_vfalu_ex1_pipex_func   (dp_vfalu_ex1_pipex_func  ),
  .dp_vfalu_ex1_pipex_imm0   (dp_vfalu_ex1_pipex_imm0  ),
  .dp_vfalu_ex1_pipex_sel    (dp_vfalu_ex1_pipex_sel   ),
  .dp_vfalu_ex1_pipex_srcf0  (dp_vfalu_ex1_pipex_srcf0 ),
  .fcnvt_ereg_forward_r_vld  (fcnvt_ereg_forward_r_vld ),
  .fcnvt_ereg_forward_result (fcnvt_ereg_forward_result),
  .fcnvt_forward_r_vld       (fcnvt_forward_r_vld      ),
  .fcnvt_forward_result      (fcnvt_forward_result     ),
  .forever_cpuclk            (forever_cpuclk           ),
  .pad_yy_icg_scan_en        (pad_yy_icg_scan_en       ),
  .vfpu_yy_xx_dqnan          (vfpu_yy_xx_dqnan         ),
  .vfpu_yy_xx_rm             (vfpu_yy_xx_rm            )
);

// &Instance("ct_fadd_top"); @28
ct_fadd_top  x_ct_fadd_top (
  .cp0_vfpu_icg_en             (cp0_vfpu_icg_en            ),
  .cp0_yy_clk_en               (cp0_yy_clk_en              ),
  .cpurst_b                    (cpurst_b                   ),
  .dp_vfalu_ex1_pipex_func     (dp_vfalu_ex1_pipex_func    ),
  .dp_vfalu_ex1_pipex_imm0     (dp_vfalu_ex1_pipex_imm0    ),
  .dp_vfalu_ex1_pipex_sel      (dp_vfalu_ex1_pipex_sel     ),
  .dp_vfalu_ex1_pipex_srcf0    (dp_vfalu_ex1_pipex_srcf0   ),
  .dp_vfalu_ex1_pipex_srcf1    (dp_vfalu_ex1_pipex_srcf1   ),
  .fadd_ereg_ex3_forward_r_vld (fadd_ereg_ex3_forward_r_vld),
  .fadd_ereg_ex3_result        (fadd_ereg_ex3_result       ),
  .fadd_forward_r_vld          (fadd_forward_r_vld         ),
  .fadd_forward_result         (fadd_forward_result        ),
  .fadd_mfvr_cmp_result        (fadd_mfvr_cmp_result       ),
  .forever_cpuclk              (forever_cpuclk             ),
  .pad_yy_icg_scan_en          (pad_yy_icg_scan_en         ),
  .vfpu_yy_xx_dqnan            (vfpu_yy_xx_dqnan           ),
  .vfpu_yy_xx_rm               (vfpu_yy_xx_rm              )
);

// &Instance("ct_fspu_top"); @29
ct_fspu_top  x_ct_fspu_top (
  .cp0_vfpu_icg_en              (cp0_vfpu_icg_en             ),
  .cp0_yy_clk_en                (cp0_yy_clk_en               ),
  .cpurst_b                     (cpurst_b                    ),
  .dp_vfalu_ex1_pipex_func      (dp_vfalu_ex1_pipex_func     ),
  .dp_vfalu_ex1_pipex_mtvr_src0 (dp_vfalu_ex1_pipex_mtvr_src0),
  .dp_vfalu_ex1_pipex_sel       (dp_vfalu_ex1_pipex_sel      ),
  .dp_vfalu_ex1_pipex_srcf0     (dp_vfalu_ex1_pipex_srcf0    ),
  .dp_vfalu_ex1_pipex_srcf1     (dp_vfalu_ex1_pipex_srcf1    ),
  .dp_vfalu_ex1_pipex_srcf2     (dp_vfalu_ex1_pipex_srcf2    ),
  .forever_cpuclk               (forever_cpuclk              ),
  .fspu_forward_r_vld           (fspu_forward_r_vld          ),
  .fspu_forward_result          (fspu_forward_result         ),
  .fspu_mfvr_data               (fspu_mfvr_data              ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          )
);

// &Instance("ct_vfalu_dp_pipe7"); @30
ct_vfalu_dp_pipe7  x_ct_vfalu_dp_pipe7 (
  .dp_vfalu_ex1_pipex_sel       (dp_vfalu_ex1_pipex_sel      ),
  .fadd_ereg_ex3_forward_r_vld  (fadd_ereg_ex3_forward_r_vld ),
  .fadd_ereg_ex3_result         (fadd_ereg_ex3_result        ),
  .fadd_forward_r_vld           (fadd_forward_r_vld          ),
  .fadd_forward_result          (fadd_forward_result         ),
  .fadd_mfvr_cmp_result         (fadd_mfvr_cmp_result        ),
  .fcnvt_ereg_forward_r_vld     (fcnvt_ereg_forward_r_vld    ),
  .fcnvt_ereg_forward_result    (fcnvt_ereg_forward_result   ),
  .fcnvt_forward_r_vld          (fcnvt_forward_r_vld         ),
  .fcnvt_forward_result         (fcnvt_forward_result        ),
  .fspu_forward_r_vld           (fspu_forward_r_vld          ),
  .fspu_forward_result          (fspu_forward_result         ),
  .fspu_mfvr_data               (fspu_mfvr_data              ),
  .pipex_dp_ex1_vfalu_mfvr_data (pipex_dp_ex1_vfalu_mfvr_data),
  .pipex_dp_ex3_vfalu_ereg_data (pipex_dp_ex3_vfalu_ereg_data),
  .pipex_dp_ex3_vfalu_freg_data (pipex_dp_ex3_vfalu_freg_data)
);


// &ModuleEnd; @32
endmodule


