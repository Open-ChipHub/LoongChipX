module slave_ram #(
    parameter int unsigned AXI_ID_WIDTH      = 7,
    parameter int unsigned AXI_ADDR_WIDTH    = 48,
    parameter int unsigned AXI_DATA_WIDTH    = 128,
    parameter int unsigned AXI_USER_WIDTH    = 2
)(
    input   logic                        clk,
    input   logic                        reset,

    input   logic                        req_i,
    input   logic                        we_i,
    input   logic [AXI_ADDR_WIDTH-1:0]   addr_i,
    input   logic [AXI_DATA_WIDTH/8-1:0] be_i,
    input   logic [AXI_DATA_WIDTH-1:0]   data_i,
    output  logic [AXI_DATA_WIDTH-1:0]   data_o
);


/// --------------------------- RAM --------------------------- ///
localparam int RamSize = 32'h400_0000 / 16;//6145;
logic [RamSize-1:0][127:0] ram_mem = {
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000030,
       128'h2e312e34_31202955_4e472820_3a434347,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_030d44d6_7000160c,
       128'h44019644_300e4400_00000044_fffff694,
       128'h000003dc_0000001c_00000000_0000030c,
       128'h44d644c1_78023016_0c440896_07814801,
       128'h800e4400_00000094_fffff62c_000003b0,
       128'h00000028_030d44d6_44c17400_160c4402,
       128'h96018148_300e4400_00000050_fffff600,
       128'h0000038c_00000020_030d44d6_44c17000,
       128'h160c4402_96018148_300e4400_0000004c,
       128'hfffff5d8_00000368_00000020_00000003,
       128'h0c44d644_c1640230_160c4408_96078148,
       128'h700e4400_00000080_fffff580_00000340,
       128'h00000024_00000003_0c44d644_c1640230,
       128'h160c4408_96078148_700e4400_00000080,
       128'hfffff528_00000318_00000024_0000030c,
       128'h44d644c1_68024016_0c440a96_09814801,
       128'h800e4400_00000084_fffff4cc_000002f0,
       128'h00000024_00030d44_d644c10e_b4030016,
       128'h0c440296_01814801_a00e4400_00000ed0,
       128'hffffe624_000002c8_00000024_00030d44,
       128'hd644c105_54030016_0c440296_01814801,
       128'ha00e4400_00000570_ffffe0dc_000002a0,
       128'h00000024_00030d44_d644c107_08030016,
       128'h0c440296_01814801_a00e4400_00000724,
       128'hffffd9e0_00000278_00000024_00030d44,
       128'hd644c101_6c030016_0c440296_01814801,
       128'ha00e4400_00000188_ffffd880_00000250,
       128'h00000024_00030d44_d644c101_6c030016,
       128'h0c440296_01814801_a00e4400_00000188,
       128'hffffd720_00000228_00000024_0000030d,
       128'h44d644c1_03340300_160c4402_96018148,
       128'h500e4400_00000350_ffffd3f8_00000200,
       128'h00000024_0000030d_44d644c1_01400300,
       128'h160c4402_96018148_600e4400_0000015c,
       128'hffffd2c4_000001d8_00000024_00000003,
       128'h0d44d644_c1740200_160c4402_96018148,
       128'h300e4400_00000090_ffffd25c_000001b0,
       128'h00000024_00000003_0d44d644_0200160c,
       128'h44019644_200e4400_00000058_ffffd228,
       128'h0000018c_00000020_00000003_0d44d654,
       128'h0200160c_44019644_300e4400_00000068,
       128'hffffd1e4_00000168_00000020_00000003,
       128'h0d44d644_c1480200_160c4402_96018148,
       128'h300e4400_00000064_ffffd1a8_00000140,
       128'h00000024_030d44d6_44c17400_160c4402,
       128'h96018148_300e4400_00000050_ffffd17c,
       128'h0000011c_00000020_030d44d6_5c00160c,
       128'h44019644_300e4400_00000030_ffffd16c,
       128'h000000fc_0000001c_030d44d6_7c00160c,
       128'h44019644_300e4400_00000050_ffffd13c,
       128'h000000dc_0000001c_030d44d6_44c16400,
       128'h160c4402_96018148_200e4400_00000040,
       128'hffffd120_000000b8_00000020_030d44d6,
       128'h44c16400_160c4402_96018148_200e4400,
       128'h00000040_ffffd104_00000094_00000020,
       128'h00000003_0d44d644_c14c0200_160c4402,
       128'h96018148_200e4400_00000068_ffffd0c4,
       128'h0000006c_00000024_00000000_00000003,
       128'h0d44d678_0200160c_44019644_300e4400,
       128'h0000008c_ffffd060_00000044_00000024,
       128'h00000000_0000030d_44d644c1_01380300,
       128'h160c4402_96018148_500e4400_00000154,
       128'hffffcf38_00000018_00000028_00030d1b,
       128'h01017801_00527a01_00000000_00000010,
       128'h412e8480_00000000_3f1a36e2_eb1c432d,
       128'h3ff00000_00000000_40180000_00000000,
       128'h40240000_00000000_402c0000_00000000,
       128'h40000000_00000000_3fe62e42_fefa39ef,
       128'h40026bb1_bbb55516_400a934f_0979a371,
       128'h3fd287a7_636f4361_3ff80000_00000000,
       128'h3fc68a28_8b60c8b3_3fd34413_509f79fb,
       128'h3fe00000_00000000_43e00000_00000000,
       128'hc1cdcd65_00000000_41cdcd65_00000000,
       128'h7fefffff_ffffffff_ffefffff_ffffffff,
       128'h41cdcd65_00000000_4197d784_00000000,
       128'h416312d0_00000000_412e8480_00000000,
       128'h40f86a00_00000000_40c38800_00000000,
       128'h408f4000_00000000_40590000_00000000,
       128'h40240000_00000000_3ff00000_00000000,
       128'hffffffff_fffff5e4_ffffffff_fffff574,
       128'hffffffff_fffff5e4_ffffffff_fffff0d8,
       128'hffffffff_fffff69c_ffffffff_fffff0d8,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffff0d8,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffff5e4_ffffffff_fffff574,
       128'hffffffff_fffff5e4_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffffa30_ffffffff_fffffa30,
       128'hffffffff_fffff9fc_ffffffff_fffff080,
       128'hffffffff_fffff09c_ffffffff_fffff09c,
       128'hffffffff_fffff09c_ffffffff_fffff09c,
       128'hffffffff_fffff09c_ffffffff_fffff048,
       128'hffffffff_fffff09c_ffffffff_fffff09c,
       128'hffffffff_fffff09c_ffffffff_fffff09c,
       128'hffffffff_fffff09c_ffffffff_fffff09c,
       128'hffffffff_fffff09c_ffffffff_ffffefb8,
       128'hffffffff_fffff09c_ffffffff_fffff064,
       128'hffffffff_fffff09c_ffffffff_fffff000,
       128'hffffffff_ffffedf0_ffffffff_ffffeea4,
       128'hffffffff_ffffeea4_ffffffff_ffffee14,
       128'hffffffff_ffffeea4_ffffffff_ffffee38,
       128'hffffffff_ffffeea4_ffffffff_ffffeea4,
       128'hffffffff_ffffeea4_ffffffff_ffffeea4,
       128'hffffffff_ffffeea4_ffffffff_ffffeea4,
       128'hffffffff_ffffeea4_ffffffff_ffffee80,
       128'hffffffff_ffffeea4_ffffffff_ffffeea4,
       128'hffffffff_ffffee5c_00000000_00696e66,
       128'h00000000_2b696e66_00000000_2d696e66,
       128'h00000000_006e616e_40140000_00000000,
       128'h40100000_00000000_40080000_00000000,
       128'h3ff00000_00000000_408f40cc_cccccccd,
       128'h00000000_00002172_65764f20_6e69614d,
       128'h00000000_00002172_6f727265_20555046,
       128'h00000000_00000a21_66252073_69202935,
       128'h642a3464_28203664_00000000_00000a21,
       128'h66252073_69203564_00000000_00000a21,
       128'h66252073_69203464_00000000_00000a21,
       128'h66252073_69203364_00000000_00000a21,
       128'h66252073_69203264_00000000_00000a21,
       128'h66252073_69203164_00000000_0000002d,
       128'h2d2d2d2d_2d2d2d55_50462074_7365542d,
       128'h2d2d2d2d_2d2d2d0a_00000000_00216d72,
       128'h6f667461_6c502068_63724167_6e6f6f4c,
       128'h206e6920_6d612049_00217364_6e656972,
       128'h46206f6c_6c65480a_4c000020_02c0c063,
       128'h28c0a076_00150184_03400000_2500018d,
       128'h28bf72cd_28ffa2cc_29ffa2cc_0320018c,
       128'h143fe20c_29bf72cc_29ff42c5_0015008c,
       128'h02c0c076_29c0a076_02ff4063_4c000020,
       128'h02c20063_28c10076_28c12061_00150184,
       128'h24ffeecc_29bfb2cc_0015008c_57eea3ff,
       128'h19fec504_001501a5_02bffc06_28fee2c7,
       128'h00150188_02ff42cd_28ff82cc_29ff62cc,
       128'h28ff02cc_29ff42cc_28ff22cc_29ff82cc,
       128'h02ff618c_28fec2cc_29fec2cc_02c0c2cc,
       128'h29c0a2cb_29c082ca_29c062c9_29c042c8,
       128'h29c022c7_29fee2c6_29ff02c5_29ff22c4,
       128'h02c14076_29c10076_29c12061_02fe0063,
       128'h4c000020_02c0c063_28c08076_28c0a061,
       128'h00150184_0015008c_57ef2fff_19fec2e4,
       128'h28ffa2c5_28ff82c6_28ff62c7_28ff42c8,
       128'h29ff42c7_29ff62c6_29ff82c5_29ffa2c4,
       128'h02c0c076_29c08076_29c0a061_02ff4063,
       128'h4c000020_02c0c063_28c08076_28c0a061,
       128'h00150184_0015008c_57ef7fff_19fec964,
       128'h00150185_02bffc06_28ff62c7_28ff42c8,
       128'h02ffa2cc_29ff42c5_29ff62c4_02c0c076,
       128'h29c08076_29c0a061_02ff4063_4c000020,
       128'h02c1c063_28c0c076_28c0e061_00150184,
       128'h24ffeecc_29bfb2cc_0015008c_57efd3ff,
       128'h19fec804_28ff62c5_28ff42c6_28ff22c7,
       128'h00150188_28ff82cc_29ff82cc_02ff618c,
       128'h28ff02cc_29ff02cc_02c0c2cc_29c0a2cb,
       128'h29c082ca_29c062c9_29c042c8_29c022c7,
       128'h29ff22c6_29ff42c5_29ff62c4_02c10076,
       128'h29c0c076_29c0e061_02fe4063_4c000020,
       128'h02c1c063_28c0c076_28c0e061_00150184,
       128'h24ffeecc_29bfb2cc_0015008c_57f053ff,
       128'h19fecc04_28ff62c5_02bffc06_28ff42c7,
       128'h00150188_28ff82cc_29ff82cc_02ff418c,
       128'h28ff22cc_29ff22cc_02c0c2cc_29c0a2cb,
       128'h29c082ca_29c062c9_29c042c8_29c022c7,
       128'h270002c6_29ff42c5_29ff62c4_02c10076,
       128'h29c0c076_29c0e061_02fe4063_4c000020,
       128'h02c20063_28c0c076_28c0e061_00150184,
       128'h24ffeecc_29bfb2cc_0015008c_57f0d3ff,
       128'h19fed404_001501a5_02bffc06_28ff22c7,
       128'h00150188_02ff62cd_28ff82cc_29ff82cc,
       128'h02ff218c_28ff02cc_29ff02cc_02c102cc,
       128'h29c0e2cb_29c0c2ca_29c0a2c9_29c082c8,
       128'h29c062c7_29c042c6_29c022c5_29ff22c4,
       128'h02c10076_29c0c076_29c0e061_02fe0063,
       128'h4c000020_02c28063_28c24076_28c26061,
       128'h00150184_0040818c_28ff62cc_4c0001a1,
       128'h00150004_28fe42c5_00150186_28fe22c7,
       128'h28fe62cd_28ff62cc_50000800_02fffd8c,
       128'h28fe22cc_680011ac_28fe22cc_28ff62cd,
       128'h47f1c19f_2800018c_28fe02cc_03400000,
       128'h29fe02cc_02c0058c_28fe02cc_4c0001a1,
       128'h001501c4_28fe42c5_00150186_28fe22c7,
       128'h28fe62cd_29ff62cd_02c0058d_28ff62cc,
       128'h2800018e_28fe02cc_50004000_29fe02cc,
       128'h02c0058c_28fe02cc_4c0001a1_02809404,
       128'h28fe42c5_00150186_28fe22c7_28fe62cd,
       128'h29ff62cd_02c0058d_28ff62cc_50007400,
       128'h29fe02cc_02c0058c_28fe02cc_29ff62c4,
       128'h57e273ff_28fe62c4_28fe42c5_28ff62c6,
       128'h28fe22c7_001501c8_00150009_0280400a,
       128'h001501ab_2700006c_24ffeacc_29c0206c,
       128'h24ffeecc_24ffe6cd_0015018e_2600018c,
       128'h29fde2cd_02c0218d_28fde2cc_50005400,
       128'h29ff62c4_57e44fff_28fe62c4_28fe42c5,
       128'h28ff62c6_28fe22c7_001501c8_00150009,
       128'h0280400a_001501ab_2700006c_24ffeacc,
       128'h29c0206c_24ffeecc_24ffe6cd_0015018e,
       128'h2600018c_29fde2cd_02c0218d_28fde2cc,
       128'h40005980_0067818c_2a3eeecc_293eeecc,
       128'h0280040c_29bfb2cc_0380858c_28bfb2cc,
       128'h29bfa2cc_0280400c_50015000_29fe02cc,
       128'h02c0058c_28fe02cc_6bffc98d_004081ad,
       128'h28bfa2cd_29bf12cd_0280058d_24ffc6cc,
       128'h4c0001a1_02808004_28fe42c5_00150186,
       128'h28fe22c7_28fe62cd_29ff62cd_02c0058d,
       128'h28ff62cc_50002800_40004580_0040818c,
       128'h0340098c_28bfb2cc_47ffa59f_29bf92cd,
       128'h02bffd8d_24ffe6cc_43ffb59f_0040818c,
       128'h0350018c_28bfb2cc_40002580_2800018c,
       128'h28ff22cc_4c0001a1_001501c4_28fe42c5,
       128'h00150186_28fe22c7_28fe62cd_29ff62cd,
       128'h02c0058d_28ff62cc_2800018e_29ff22cd,
       128'h02c0058d_28ff22cc_50003800_6bffc98d,
       128'h004081ad_28bfa2cd_29bf12cd_0280058d,
       128'h24ffc6cc_4c0001a1_02808004_28fe42c5,
       128'h00150186_28fe22c7_28fe62cd_29ff62cd,
       128'h02c0058d_28ff62cc_50002800_44007d80,
       128'h0040818c_0340098c_28bfb2cc_29bf12cc,
       128'h001531ac_001331cc_0013b1ad_004081ed,
       128'h0012b58c_0040818c_0040818e_004081ad,
       128'h28bf92cf_28bf92cd_28bf12cc_40003580,
       128'h0040818c_0350018c_28bfb2cc_29bf12cc,
       128'h0015008c_57de9bff_28ff22c4_00150185,
       128'h02bffc0c_50000800_2abf92cc_40000d80,
       128'h0040818c_28bf92cc_29ff22cc_2600018c,
       128'h29fde2cd_02c0218d_28fde2cc_5002e400,
       128'h29fe02cc_02c0058c_28fe02cc_6bffc98d,
       128'h004081ad_28bfa2cd_29bf42cd_0280058d,
       128'h24ffd2cc_4c0001a1_02808004_28fe42c5,
       128'h00150186_28fe22c7_28fe62cd_29ff62cd,
       128'h02c0058d_28ff62cc_50002800_40004580,
       128'h0040818c_0340098c_28bfb2cc_4c0001a1,
       128'h001501c4_28fe42c5_00150186_28fe22c7,
       128'h28fe62cd_29ff62cd_02c0058d_28ff62cc,
       128'h00005d8e_2400018c_29fde2cd_02c0218d,
       128'h28fde2cc_6bffc98d_004081ad_28bfa2cd,
       128'h29bf42cd_0280058d_24ffd2cc_4c0001a1,
       128'h02808004_28fe42c5_00150186_28fe22c7,
       128'h28fe62cd_29ff62cd_02c0058d_28ff62cc,
       128'h50002800_44004580_0040818c_0340098c,
       128'h28bfb2cc_29bf42cc_0280040c_5003d400,
       128'h29fe02cc_02c0058c_28fe02cc_29ff62c4,
       128'h57f007ff_28fe62c4_28fe42c5_28ff62c6,
       128'h28fe22c7_00150188_001501a9_001501ca,
       128'h24ffe6cc_24ffeacd_24ffeece_2b800180,
       128'h29fde2cd_02c0218d_28fde2cc_29bfb2cc,
       128'h0380818c_28bfb2cc_5c0011ac_02811c0c,
       128'h0015018d_2800018c_28fe02cc_580019ac,
       128'h0281140c_0015018d_2800018c_28fe02cc,
       128'h29bfb2cc_03a0018c_28bfb2cc_5c0011ac,
       128'h02811c0c_0015018d_2800018c_28fe02cc,
       128'h580019ac_02819c0c_0015018d_2800018c,
       128'h28fe02cc_50048c00_29fe02cc_02c0058c,
       128'h28fe02cc_29ff62c4_57e99bff_28fe62c4,
       128'h28fe42c5_28ff62c6_28fe22c7_00150188,
       128'h001501a9_001501ca_24ffe6cc_24ffeacd,
       128'h24ffeece_2b800180_29fde2cd_02c0218d,
       128'h28fde2cc_29bfb2cc_0380818c_28bfb2cc,
       128'h5c0011ac_0281180c_0015018d_2800018c,
       128'h28fe02cc_5004fc00_29fe02cc_02c0058c,
       128'h28fe02cc_29ff62c4_57e6fbff_28fe62c4,
       128'h28fe42c5_28ff62c6_28fe22c7_001501a8,
       128'h00150009_001501ca_001501eb_2700006c,
       128'h24ffeacc_29c0206c_24ffeecc_24ffe6cf,
       128'h2abf52ce_2abed2cd_29bed2cc_2400018c,
       128'h29fde2cd_02c0218d_28fde2cc_50001400,
       128'h0040818c_006f818c_2400018c_29fde2cd,
       128'h02c0218d_28fde2cc_40002180_0040818c,
       128'h0342018c_28bfb2cc_50004000_0040818c,
       128'h0067818c_2400018c_29fde2cd_02c0218d,
       128'h28fde2cc_40002180_0040818c_0341018c,
       128'h28bfb2cc_5000b400_29ff62c4_57e7afff,
       128'h28fe62c4_28fe42c5_28ff62c6_28fe22c7,
       128'h001501a8_00150009_001501ca_001501eb,
       128'h2700006c_24ffeacc_29c0206c_24ffeecc,
       128'h24ffe6cf_2abf52ce_2600018d_29fde2cd,
       128'h02c0218d_28fde2cc_40005980_0040818c,
       128'h0344018c_28bfb2cc_50011800_29ff62c4,
       128'h57e99bff_28fe62c4_28fe42c5_28ff62c6,
       128'h28fe22c7_001501a8_00150009_001501ca,
       128'h001501eb_2700006c_24ffeacc_29c0206c,
       128'h24ffeecc_24ffe6cf_2abf52ce_2600018d,
       128'h29fde2cd_02c0218d_28fde2cc_40005980,
       128'h0040818c_0348018c_28bfb2cc_50017c00,
       128'h29ff62c4_57e877ff_28fe62c4_28fe42c5,
       128'h28ff62c6_28fe22c7_001501a8_001501c9,
       128'h001501ea_0015020b_2700006c_24ffeacc,
       128'h29c0206c_24ffeecc_24ffe6d0_2abf52cf,
       128'h0067818e_0044fd8c_28bec2cc_00df018d,
       128'h0040818c_001131ac_0015b58d_28bec2cd,
       128'h0048fd8c_28bec2cc_29bec2cc_2400018c,
       128'h29fde2cd_02c0218d_28fde2cc_50001400,
       128'h0000598c_2400018c_29fde2cd_02c0218d,
       128'h28fde2cc_40001d80_0040818c_0342018c,
       128'h28bfb2cc_50003c00_00005d8c_2400018c,
       128'h29fde2cd_02c0218d_28fde2cc_40001d80,
       128'h0040818c_0341018c_28bfb2cc_50024c00,
       128'h29ff62c4_57e947ff_28fe62c4_28fe42c5,
       128'h28ff62c6_28fe22c7_00150208_001501a9,
       128'h001501ca_001501eb_2700006c_24ffeacc,
       128'h29c0206c_24ffeecc_24ffe6cf_2abf52ce,
       128'h0067818d_0045fd8c_28fea2cc_00150190,
       128'h0011b58c_0015b1ac_28fea2cc_0049fd8d,
       128'h28fea2cc_29fea2cc_2600018c_29fde2cd,
       128'h02c0218d_28fde2cc_40008180_0040818c,
       128'h0344018c_28bfb2cc_5002d800_29ff62c4,
       128'h57eb5bff_28fe62c4_28fe42c5_28ff62c6,
       128'h28fe22c7_00150208_001501a9_001501ca,
       128'h001501eb_2700006c_24ffeacc_29c0206c,
       128'h24ffeecc_24ffe6cf_2abf52ce_0067818d,
       128'h0045fd8c_28fe82cc_00150190_0011b58c,
       128'h0015b1ac_28fe82cc_0049fd8d_28fe82cc,
       128'h29fe82cc_2600018c_29fde2cd_02c0218d,
       128'h28fde2cc_40008180_0040818c_0348018c,
       128'h28bfb2cc_5c01edac_0281900c_0015018d,
       128'h2800018c_28fe02cc_580019ac_0281a40c,
       128'h0015018d_2800018c_28fe02cc_29bfb2cc,
       128'h0014b1ac_02bff80c_28bfb2cd_40001580,
       128'h0040818c_0350018c_28bfb2cc_29bfb2cc,
       128'h0014b1ac_02bfcc0c_28bfb2cd_580015ac,
       128'h0281900c_0015018d_2800018c_28fe02cc,
       128'h580029ac_0281a40c_0015018d_2800018c,
       128'h28fe02cc_29bfb2cc_0380818c_28bfb2cc,
       128'h5c0011ac_0281600c_0015018d_2800018c,
       128'h28fe02cc_29bfb2cc_0014b1ac_02bfbc0c,
       128'h28bfb2cd_29bf52cc_0280280c_50001c00,
       128'h29bf52cc_0280080c_5c0011ac_0281880c,
       128'h0015018d_2800018c_28fe02cc_50003c00,
       128'h29bf52cc_0280200c_5c0011ac_0281bc0c,
       128'h0015018d_2800018c_28fe02cc_50005c00,
       128'h29bf52cc_0280400c_5c0011ac_0281600c,
       128'h0015018d_2800018c_28fe02cc_580019ac,
       128'h0281e00c_0015018d_2800018c_28fe02cc,
       128'h50095c00_67ff6dcd_0281a40d_0015018e,
       128'h60096dae_0281e00d_0015018e_4c000180,
       128'h0010b1ac_18007a8c_2600018d_0010b1ac,
       128'h18007aec_00410d8d_00df01cc_6809998d,
       128'h0281080c_004081cd_0015018e_02bf6d8c,
       128'h5009ac00_44070d80_0067818c_0012b00c,
       128'h0350018c_4408b1a0_006781ad_0012b40d,
       128'h0342018d_440079a0_006781ad_0012b40d,
       128'h0014b58d_038105ad_1400012d_0018b1ac,
       128'h0280040d_0040818c_02be5d8c_5009f800,
       128'h640055cd_0280940d_0015018e_600095ae,
       128'h02819c0d_0015018e_2800018c_28fe02cc,
       128'h03400000_50000800_03400000_50001000,
       128'h03400000_50001800_29fe02cc_02c0058c,
       128'h28fe02cc_29bfb2cc_0384018c_28bfb2cc,
       128'h50003400_29fe02cc_02c0058c_28fe02cc,
       128'h29bfb2cc_0384018c_28bfb2cc_50005000,
       128'h29fe02cc_02c0058c_28fe02cc_29bfb2cc,
       128'h0384018c_28bfb2cc_50006800_29fe02cc,
       128'h02c0058c_28fe02cc_29bfb2cc_0381018c,
       128'h28bfb2cc_5c0085ac_0281a00c_0015018d,
       128'h2800018c_28fe02cc_29fe02cc_02c0058c,
       128'h28fe02cc_29bfb2cc_0382018c_28bfb2cc,
       128'h5000a800_29fe02cc_02c0058c_28fe02cc,
       128'h29bfb2cc_0388018c_28bfb2cc_5c00c5ac,
       128'h0281b00c_0015018d_2800018c_28fe02cc,
       128'h29fe02cc_02c0058c_28fe02cc_29bfb2cc,
       128'h0384018c_28bfb2cc_4c000180_0010b1ac,
       128'h180082ac_2600018d_0010b1ac_1800830c,
       128'h00410d8d_00df01cc_6801098d_0280480c,
       128'h004081cd_0015018e_02be618c_2800018c,
       128'h28fe02cc_29fe02cc_02c0058c_28fe02cc,
       128'h29bf92cc_0040818c_0013b58c_020001ad,
       128'h004081ad_28bef2cc_28bef2cd_29bef2cc,
       128'h2400018c_29fde2cd_02c0218d_28fde2cc,
       128'h5c0041ac_0280a80c_0015018d_2800018c,
       128'h28fe02cc_50005400_29bf92cc_0015008c,
       128'h57e897ff_00150184_02fe02cc_40001d80,
       128'h0015008c_57e853ff_00150184_2800018c,
       128'h28fe02cc_29fe02cc_02c0058c_28fe02cc,
       128'h29bfb2cc_0390018c_28bfb2cc_5c009dac,
       128'h0280b80c_0015018d_2800018c_28fe02cc,
       128'h29bf92c0_29fe02cc_02c0058c_28fe02cc,
       128'h29bfa2cc_28bf02cc_50000c00_29bfa2cc,
       128'h0040818c_0011300c_28bf02cc_29bfb2cc,
       128'h0380098c_28bfb2cc_64002580_0040818c,
       128'h28bf02cc_29bf02cc_2400018c_29fde2cd,
       128'h02c0218d_28fde2cc_5c0059ac_0280a80c,
       128'h0015018d_2800018c_28fe02cc_50006c00,
       128'h29bfa2cc_0015008c_57e95fff_00150184,
       128'h02fe02cc_40001d80_0015008c_57e91bff,
       128'h00150184_2800018c_28fe02cc_29bfa2c0,
       128'h47ff019f_0040818c_28bf82cc_03400000,
       128'h29bf82c0_50000c00_29bf82cc_0280040c,
       128'h29fe02cc_02c0058c_28fe02cc_29bfb2cc,
       128'h0380418c_28bfb2cc_50003000_29bf82cc,
       128'h0280040c_29fe02cc_02c0058c_28fe02cc,
       128'h29bfb2cc_0380218c_28bfb2cc_50005400,
       128'h29bf82cc_0280040c_29fe02cc_02c0058c,
       128'h28fe02cc_29bfb2cc_0380118c_28bfb2cc,
       128'h50007800_29bf82cc_0280040c_29fe02cc,
       128'h02c0058c_28fe02cc_29bfb2cc_0380098c,
       128'h28bfb2cc_50009c00_29bf82cc_0280040c,
       128'h29fe02cc_02c0058c_28fe02cc_29bfb2cc,
       128'h0380058c_28bfb2cc_4c000180_0010b1ac,
       128'h180090ec_2600018d_0010b1ac_1800914c,
       128'h00410d8d_00df01cc_6800d98d_0280400c,
       128'h004081cd_0015018e_02bf818c_2800018c,
       128'h28fe02cc_29bfb2c0_29fe02cc_02c0058c,
       128'h28fe02cc_500dec00_29fe02cc_02c0058c,
       128'h28fe02cc_4c0001a1_001501c4_28fe42c5,
       128'h00150186_28fe22c7_28fe62cd_29ff62cd,
       128'h02c0058d_28ff62cc_2800018e_28fe02cc,
       128'h580041ac_0280940c_0015018d_2800018c,
       128'h28fe02cc_500e3c00_29fe62cc_19ff4a6c,
       128'h440e4980_28fe42cc_29ff62c0_29fde2c8,
       128'h29fe02c7_29fe22c6_29fe42c5_29fe62c4,
       128'h02c28076_29c24076_29c26061_02fd8063,
       128'h4c000020_02c28063_28c24076_28c26061,
       128'h00150184_28fe62cc_6bffcdac_2abe02cc,
       128'h0011b1ad_28ff02cc_28fe62cd_4c0001a1,
       128'h02808004_28fe82c5_00150186_28fe42c7,
       128'h28fea2cd_29fe62cd_02c0058d_28fe62cc,
       128'h50002800_40004180_0040818c_0340098c,
       128'h28bdf2cc_29fe62c4_57f0cbff_28fea2c4,
       128'h28fe82c5_28fe62c6_28fe42c7_001501e8,
       128'h001501c9_0280280a_0015000b_2700006c,
       128'h29c0206d_0280140d_0040818c_02bffd8c,
       128'h28bfa2cc_0067818e_0044fd8c_28bfb2cc,
       128'h0015018f_0040818c_001131ac_0015b58d,
       128'h28bfb2cd_0048fd8c_28bfb2cc_4c0001c1,
       128'h00150184_28fe82c5_001501a6_28fe42c7,
       128'h28fea2ce_29fe62ce_02c005ae_28fe62cd,
       128'h0281940c_50000800_0281140c_40000d80,
       128'h0040818c_0340818c_28bdf2cc_4000f980,
       128'h0040818c_28bfa2cc_29fe62c4_57f48fff,
       128'h28fea2c4_28fe82c5_28fe62c6_28fe42c7,
       128'h00150188_001501a9_001501ca_24ff86cc,
       128'h24ffe6cd_0040818e_0014b1ac_039ffd8c,
       128'h15ffffec_28bdf2cd_2bbe22c0_50000800,
       128'h01141800_2bbe22c0_40001180_0067818c,
       128'h2a3f8ecc_29ff02cc_28fe62cc_2bfe22c0,
       128'h01070020_2bbe22c1_2bbee2c0_40001580,
       128'h0040818c_28bfb2cc_29bf92c0_40000980,
       128'h0040818c_28bfa2cc_40001580_0040818c,
       128'h0340098c_28bdf2cc_29bf92c0_50000800,
       128'h29bf92cc_001131ac_28bfa2cc_28bf92cd,
       128'h6c00198d_0040818c_004081ad_28bfa2cc,
       128'h28be02cd_29bf92cc_28be02cc_29be12cc,
       128'h02bffd8c_28be12cc_40001180_0040818c,
       128'h0350018c_28bdf2cc_40002180_0040818c,
       128'h28be12cc_50002c00_29bfb2c0_29bfa2c0,
       128'h29bdf2cc_0390018c_28bdf2cc_29be12c0,
       128'h50000800_29be12cc_0040818c_02bffd8c,
       128'h0040818c_001131ac_28bfb2cc_24ff86cd,
       128'h6400258d_0040818c_28bfb2cc_24ff86cd,
       128'h48005000_0c218020_2b800180_1800cbcc,
       128'h2bbe22c1_48006400_0c238400_2b800180,
       128'h1800cc2c_2bbe22c1_4000a180_0040818c,
       128'h0360018c_28bdf2cc_29bfa2cc_0280140c,
       128'h50000800_0280100c_60000dac_02be740c,
       128'h0040818d_28bfb2cc_60001d8d_02818c0c,
       128'h0040818d_28bfb2cc_2bfee2c0_01070020,
       128'h2b800180_1800ce0c_2bbee2c1_29bfb2cc,
       128'h02bffd8c_28bfb2cc_48002400_0c218020,
       128'h2bbe22c1_2bbee2c0_2bfee2c0_01050020,
       128'h01010040_2b800180_1800d02c_01070042,
       128'h01010060_01070080_2bbf22c4_01010080,
       128'h2b800180_1800d0cc_01070084_2bbf22c4,
       128'h01010080_2b800180_1800d12c_01070084,
       128'h2b800180_1800d14c_2bbf22c4_01030063,
       128'h2bbf42c0_2b800183_1800d1ac_01010002,
       128'h2bbf42c0_2bbee2c1_29fee2cc_0041d18c,
       128'h0040818c_028ffd8c_28bf72cc_2bff22c0,
       128'h01050000_2bbf42c0_2bff42c0_01030020,
       128'h01050040_2b800180_1800d36c_011d2002,
       128'h2b3f72c0_01050021_2b800180_1800d3cc,
       128'h011d2001_2b3fb2c0_29bf72cc_0114b40c,
       128'h011a8800_01010020_2b800180_1800d34c,
       128'h01050021_2b800180_1800d4ec_011d2001,
       128'h2b3fb2c0_29bfb2cc_0114b40c_011a8800,
       128'h01010020_01050040_2b800180_1800d5cc,
       128'h01030042_2b800180_1800d5ec_2bbee2c2,
       128'h01010021_2b800180_1800d62c_01050021,
       128'h2b800180_1800d64c_011d2001_2b3f72c0,
       128'h29fee2cc_001531ac_030ffd8c_0015000c,
       128'h0014b1ad_0300018c_02bffc0c_28fee2cd,
       128'h29bf72cc_02b0058c_0040818c_035ffd8c,
       128'h0040818c_0045d18c_28fee2cc_2bfee2c0,
       128'h2bbe22c0_29be12cc_0280180c_44000d80,
       128'h0040818c_0350018c_28bdf2cc_2bfe22c0,
       128'h01141800_2bbe22c0_40001180_0067818c,
       128'h2a3f8ecc_293f8ecc_0114b40c_0114d400,
       128'h0c218400_0114a801_2bbe22c0_5004ac00,
       128'h0015008c_57f837ff_28fea2c4_28fe82c5,
       128'h28fe62c6_28fe42c7_2bbe22c0_00150188,
       128'h001501a9_001501ca_24ff86cc_24ff82cd,
       128'h24ff7ece_48003c00_0c218020_2b800180,
       128'h1800dbac_2bbe22c1_48001900_0c218400,
       128'h2b800180_1800dc8c_2bbe22c1_48002d00,
       128'h0c2c0020_2bbe22c0_2bbe22c1_29bdf2cc,
       128'h001501ac_29be02cc_001501cc_29be12cc,
       128'h0015014d_0015012e_0015010c_2bfe22c0,
       128'h29fe42c7_29fe62c6_29fe82c5_29fea2c4,
       128'h02c28076_29c24076_29c26061_02fd8063,
       128'h4c000020_02c28063_28c24076_28c26061,
       128'h00150184_0015008c_57f13fff_28fe62c4,
       128'h28fe42c5_28fe22c6_28fe02c7_001501c8,
       128'h28ffa2c9_0015018a_001501ab_02fe82ce,
       128'h24ff72cc_24ff6ecd_293ec1ac_0280800c,
       128'h0010d98d_02ffc18c_29ffa2cd_02c0058d,
       128'h28ffa2cc_40002180_0040818c_0340218c,
       128'h28bdb2cc_50003000_293ec1ac_0280ac0c,
       128'h0010d98d_02ffc18c_29ffa2cd_02c0058d,
       128'h28ffa2cc_40002580_0040818c_0340118c,
       128'h28bdb2cc_50006000_293ec1ac_0280b40c,
       128'h0010d98d_02ffc18c_29ffa2cd_02c0058d,
       128'h28ffa2cc_40002580_0067818c_2a3f9ecc,
       128'h68008d8d_02807c0c_28ffa2cd_6fffd18d,
       128'h02807c0c_28ffa2cd_6c0011ac_28ffa2cd,
       128'h2abdc2cc_293ec1ac_0280c00c_0010d98d,
       128'h02ffc18c_29ffa2cd_02c0058d_28ffa2cc,
       128'h50002000_29bdc2cc_02bffd8c_28bdc2cc,
       128'h40003180_0040818c_0340318c_28bdb2cc,
       128'h44001580_0067818c_2a3f9ecc_40004d80,
       128'h0040818c_28bdc2cc_40007180_0040818c,
       128'h0340058c_28bdb2cc_44008180_0040818c,
       128'h0340098c_28bdb2cc_03400000_50000800,
       128'h6fff7d8d_02807c0c_28ffa2cd_40001580,
       128'h0040818c_28bf82cc_29bf82cc_001501ac,
       128'h002a0007_5c000980_002031ad_0040818c,
       128'h004081ad_0280280c_28bf82cd_293ec1ac,
       128'h0010d9ad_02ffc1ad_00005dcc_29ffa2cc,
       128'h02c005ac_28ffa2cd_0067818e_0280c18c,
       128'h0067818c_0040818c_001501ac_002a0007,
       128'h5c000980_0020b1ad_0040818c_004081ad,
       128'h0280280c_28bf82cd_50008000_293ec1ac,
       128'h0280b80c_0010d98d_02ffc18c_29ffa2cd,
       128'h02c0058d_28ffa2cc_6800a18d_02807c0c,
       128'h28ffa2cd_47ffcd9f_29bf52cd_02bffd8d,
       128'h24ffd6cc_6800158d_02807c0c_28ffa2cd,
       128'h293ec1ac_0280c00c_0010d98d_02ffc18c,
       128'h29ffa2cd_02c0058d_28ffa2cc_50002000,
       128'h03400000_50002800_6fff918d_02807c0c,
       128'h28ffa2cd_40001580_28ff62cc_29ff62cc,
       128'h002a0007_5c0009a0_0023358c_0280280d,
       128'h28ff62cc_293ec1ac_0010d9ad_02ffc1ad,
       128'h00005dcc_29ffa2cc_02c005ac_28ffa2cd,
       128'h0067818e_0280c18c_006781ac_002a0007,
       128'h5c000980_0023b1ad_0280280c_28ff62cd,
       128'h29bf52cc_02bffd8c_28bf52cc_50006c00,
       128'h29bf52cc_28bdd2cc_50017000_29bf82cc,
       128'h0280058c_28bf82cc_40018180_0040818c,
       128'h0340058c_28bf82cc_48011000_0c218400,
       128'h2b800180_1800f90c_2bbf22c1_44001980,
       128'h0067818c_03c0058c_0067818c_0114b40c,
       128'h0114d400_0c218020_2b800180_1800fa4c,
       128'h2bbf22c1_2bff22c0_01030020_2bbde2c1,
       128'h011d2000_2b3f82c0_44007580_0040818c,
       128'h28bdd2cc_29ff62cc_02c0058c_28ff62cc,
       128'h40001180_0340058c_28ff62cc_40001180,
       128'h28ff62cc_48002500_0c218020_2b800180,
       128'h1800fcec_2bbf22c1_50003800_29bf82cc,
       128'h0280058c_28bf82cc_29ff62c0_48004c00,
       128'h0c238020_2b800181_0010b1ac_00410d8c,
       128'h2abdd2cc_1800facd_01010000_011d2800,
       128'h0114a980_0015358c_004505ad_28ff62cd,
       128'h0340058c_28ff62cc_50002400_011d2800,
       128'h0114a980_28ff62cc_60001580_28ff62cc,
       128'h29ff62cc_02c0058c_28ff62cc_48007800,
       128'h0c218400_2b800180_1801012c_2bbf22c1,
       128'h2bff22c0_01030020_2bbf02c1_01010000,
       128'h011d2800_0114a980_0015358c_004505ad,
       128'h28ff62cd_0340058c_28ff62cc_50002400,
       128'h011d2800_0114a980_28ff62cc_60001580,
       128'h28ff62cc_29ff62cd_001531ad_0114b80d,
       128'h011aa800_0041818c_1600000c_1500000c,
       128'h01030400_50002000_0114b80d_011aa800,
       128'h48001100_0c238020_2b800181_1801050c,
       128'h2bbf02c0_2bff02c0_01050020_2b800180,
       128'h0010b1ac_00410d8c_2abdd2cc_1801028d,
       128'h01030021_2bbde2c1_011d2000_2b3f82c0,
       128'h29bf82cc_0114b40c_011a8800_2bbde2c0,
       128'h6bffc18d_0280240c_0040818d_28bdd2cc,
       128'h6800158d_02807c0c_28ffa2cd_29bdd2cc,
       128'h02bffd8c_28bdd2cc_293ec1ac_0280c00c,
       128'h0010d98d_02ffc18c_29ffa2cd_02c0058d,
       128'h28ffa2cc_50002c00_29bdd2cc_0280180c,
       128'h44003980_0040818c_0350018c_28bdb2cc,
       128'h2bfde2c0_01030020_2bbde2c0_0114a801,
       128'h293f9ecc_0280040c_48001c00_0c218400,
       128'h0114a801_2bbde2c0_293f9ec0_50055c00,
       128'h0015008c_54057800_28fe62c4_28fe42c5,
       128'h28fe22c6_28fe02c7_2bbde2c0_00150188,
       128'h001501a9_001501ca_24ff76cc_24ff72cd,
       128'h24ff6ece_48003c00_0c218020_2b800180,
       128'h18010d6c_2bbde2c1_48001900_0c218400,
       128'h2b800180_18010dcc_2bbde2c1_5005bc00,
       128'h0015008c_57f6fbff_28fe62c4_28fe42c5,
       128'h28fe22c6_28fe02c7_00150188_001501a9,
       128'h001501ca_001501eb_24ff72ce_24ff6ecf,
       128'h02800c0d_50000800_0280100d_40000da0,
       128'h004081ad_034011ad_28bdb2cd_1800f38c,
       128'h50000800_1800f38c_40000d80_0040818c,
       128'h0340118c_28bdb2cc_48007000_0c218400,
       128'h2b800180_1801118c_2bbde2c1_50063c00,
       128'h0015008c_57f77bff_28fe62c4_28fe42c5,
       128'h28fe22c6_28fe02c7_1800f568_02801009,
       128'h0015018a_001501ab_24ff72cc_24ff6ecd,
       128'h48003800_0c218020_2b800180_1801138c,
       128'h2bbde2c1_50068400_0015008c_57f7c3ff,
       128'h28fe62c4_28fe42c5_28fe22c6_28fe02c7,
       128'h1800f768_02800c09_0015018a_001501ab,
       128'h24ff72cc_24ff6ecd_48003900_0c220020,
       128'h2bbde2c0_2bbde2c1_29ff22c0_29ffa2c0,
       128'h29bdb2cc_001501ac_29bdc2cc_001501cc,
       128'h29bdd2cc_0015014d_0015012e_0015010c,
       128'h2bfde2c0_29fe02c7_29fe22c6_29fe42c5,
       128'h29fe62c4_02c28076_29c24076_29c26061,
       128'h02fd8063_4c000020_02c28063_28c24076,
       128'h28c26061_00150184_0015008c_57f9bfff,
       128'h28fee2c4_28fec2c5_28fea2c6_28fe82c7,
       128'h001501e8_28ffa2c9_001501aa_001501cb,
       128'h2700006c_24ff92cc_29c0206c_240002cc,
       128'h29c0406c_24000acc_02ff02cf_2a3e5ecd,
       128'h0040818e_28fe22cc_6fff518d_02807c0c,
       128'h28ffa2cd_40001180_28fe62cc_29fe62cc,
       128'h002a0007_5c0009a0_0023358c_28fe22cd,
       128'h28fe62cc_293f41ac_0010d9ad_02ffc1ad,
       128'h29ffa2ce_02c005ae_28ffa2cd_00005d8c,
       128'h0067818c_02bfd98c_0067818c_0010358c,
       128'h2a3f9ecd_0281840c_50000800_0281040c,
       128'h40000d80_0040818c_0340818c_288022cc,
       128'h50003800_00005d8c_0067818c_0280c18c,
       128'h2a3f9ecc_6000198d_0280240c_00005d8d,
       128'h2a3f9ecc_293f9ecc_002a0007_5c0009a0,
       128'h0023b58c_28fe22cd_28fe62cc_4000b980,
       128'h28fe62cc_40000d80_0040818c_0350018c,
       128'h288022cc_298022cc_0014b1ac_02bfbc0c,
       128'h288022cd_44001580_28fe62cc_29ffa2c0,
       128'h29be42cc_001501ac_293e5ecc_0015016d,
       128'h29fe22ca_0015012c_29fe62c8_29fe82c7,
       128'h29fea2c6_29fec2c5_29fee2c4_02c28076,
       128'h29c24076_29c26061_02fd8063_4c000020,
       128'h02c28063_28c24076_28c26061_00150184,
       128'h0015008c_57fb47ff_28fee2c4_28fec2c5,
       128'h28fea2c6_28fe82c7_001501e8_28ffa2c9,
       128'h001501aa_001501cb_2700006c_24ff92cc,
       128'h29c0206c_240002cc_29c0406c_24000acc,
       128'h02ff02cf_2a3e5ecd_0040818e_28fe22cc,
       128'h6fff518d_02807c0c_28ffa2cd_40001180,
       128'h28fe62cc_29fe62cc_002a0007_5c0009a0,
       128'h0023358c_28fe22cd_28fe62cc_293f41ac,
       128'h0010d9ad_02ffc1ad_29ffa2ce_02c005ae,
       128'h28ffa2cd_00005d8c_0067818c_02bfd98c,
       128'h0067818c_0010358c_2a3f9ecd_0281840c,
       128'h50000800_0281040c_40000d80_0040818c,
       128'h0340818c_288022cc_50003800_00005d8c,
       128'h0067818c_0280c18c_2a3f9ecc_6000198d,
       128'h0280240c_00005d8d_2a3f9ecc_293f9ecc,
       128'h002a0007_5c0009a0_0023b58c_28fe22cd,
       128'h28fe62cc_4000b980_28fe62cc_40000d80,
       128'h0040818c_0350018c_288022cc_298022cc,
       128'h0014b1ac_02bfbc0c_288022cd_44001580,
       128'h28fe62cc_29ffa2c0_29be42cc_001501ac,
       128'h293e5ecc_0015016d_29fe22ca_0015012c,
       128'h29fe62c8_29fe82c7_29fea2c6_29fec2c5,
       128'h29fee2c4_02c28076_29c24076_29c26061,
       128'h02fd8063_4c000020_02c14063_28c10076,
       128'h28c12061_00150184_0015008c_57fb73ff,
       128'h28ffa2c4_28ff82c5_28ff62c6_28ff42c7,
       128'h28ff22c8_28ff02c9_0015018a_001501ab,
       128'h24000acc_240012cd_2900018d_0280800d,
       128'h0010b1ac_28ff22cd_29ff02cd_02c0058d,
       128'h28ff02cc_40002180_0040818c_0340218c,
       128'h288042cc_50003000_2900018d_0280ac0d,
       128'h0010b1ac_28ff22cd_29ff02cd_02c0058d,
       128'h28ff02cc_40002580_0040818c_0340118c,
       128'h288042cc_50006000_2900018d_0280b40d,
       128'h0010b1ac_28ff22cd_29ff02cd_02c0058d,
       128'h28ff02cc_40002580_0067818c_2a3efecc,
       128'h68008d8d_02807c0c_28ff02cd_2900018d,
       128'h0280c00d_0010b1ac_28ff22cd_29ff02cd,
       128'h02c0058d_28ff02cc_6800218d_02807c0c,
       128'h28ff02cd_2900018d_0281880d_0010b1ac,
       128'h28ff22cd_29ff02cd_02c0058d_28ff02cc,
       128'h6800218d_02807c0c_28ff02cd_5c002dac,
       128'h0280080c_0040818d_28bee2cc_50003c00,
       128'h2900018d_0281600d_0010b1ac_28ff22cd,
       128'h29ff02cd_02c0058d_28ff02cc_6800258d,
       128'h02807c0c_28ff02cd_40003180_0040818c,
       128'h0340818c_288042cc_5c0041ac_0280400c,
       128'h0040818d_28bee2cc_50008800_2900018d,
       128'h0281e00d_0010b1ac_28ff22cd_29ff02cd,
       128'h02c0058d_28ff02cc_6800258d_02807c0c,
       128'h28ff02cd_44003180_0040818c_0340818c,
       128'h288042cc_5c0041ac_0280400c_0040818d,
       128'h28bee2cc_29ff02cc_02fffd8c_28ff02cc,
       128'h5c0011ac_0280400c_0040818d_28bee2cc,
       128'h40002180_28ff02cc_29ff02cc_02fffd8c,
       128'h28ff02cc_5c0035ac_28ff02cd_2a8022cc,
       128'h580011ac_28ff02cd_2a8002cc_40004d80,
       128'h28ff02cc_44005580_0040818c_0350018c,
       128'h288042cc_40015d80_0040818c_0340418c,
       128'h288042cc_6fffc18d_02807c0c_28ff02cd,
       128'h6c0011ac_28ff02cd_2a8022cc_40001d80,
       128'h0040818c_0340058c_288042cc_2900018d,
       128'h0280c00d_0010b1ac_28ff22cd_29ff02cd,
       128'h02c0058d_28ff02cc_50002000_6fffd18d,
       128'h02807c0c_28ff02cd_6c0031ac_28ff02cd,
       128'h2a8002cc_2900018d_0280c00d_0010b1ac,
       128'h28ff22cd_29ff02cd_02c0058d_28ff02cc,
       128'h50002000_298022cc_02bffd8c_288022cc,
       128'h40003180_0040818c_0340318c_288042cc,
       128'h44001580_0067818c_2a3efecc_40004d80,
       128'h0040818c_0340058c_288042cc_40005d80,
       128'h0040818c_288022cc_4400c980_0040818c,
       128'h0340098c_288042cc_29bee2cc_001501ac,
       128'h293efecc_0015016d_0015014c_29ff02c9,
       128'h29ff22c8_29ff42c7_29ff62c6_29ff82c5,
       128'h29ffa2c4_02c14076_29c10076_29c12061,
       128'h02fec063_4c000020_02c18063_28c14076,
       128'h28c16061_00150184_28ff22cc_6bffcdac,
       128'h2abeb2cc_0011b1ad_28ff82cc_28ff22cd,
       128'h4c0001a1_02808004_28ff42c5_00150186,
       128'h28ff02c7_28ff62cd_29ff22cd_02c0058d,
       128'h28ff22cc_50002800_40004180_0040818c,
       128'h0340098c_28bea2cc_47ffbd9f_28fec2cc,
       128'h4c0001a1_001501c4_28ff42c5_00150186,
       128'h28ff02c7_28ff62cd_29ff22cd_02c0058d,
       128'h28ff22cc_2800018e_0010b1ac_28fec2cc,
       128'h28fee2cd_29fec2cc_02fffd8c_28fec2cc,
       128'h50004400_6bffc9ac_28ffa2cd_2abeb2cc,
       128'h29ffa2cc_02c0058c_28ffa2cc_4c0001a1,
       128'h02808004_28ff42c5_00150186_28ff02c7,
       128'h28ff62cd_29ff22cd_02c0058d_28ff22cc,
       128'h50003400_29ffa2cc_28fec2cc_44009180,
       128'h0040818c_0340058c_28bea2cc_4400a180,
       128'h0040818c_0340098c_28bea2cc_29ff82cc,
       128'h28ff22cc_29bea2cc_001501ac_29beb2cc,
       128'h0015016d_0015014c_29fec2c9_29fee2c8,
       128'h29ff02c7_29ff22c6_29ff42c5_29ff62c4,
       128'h02c18076_29c14076_29c16061_02fe8063,
       128'h4c000020_02c0c063_28c08076_28c0a061,
       128'h00150184_24ffeecc_47ffa99f_0015008c,
       128'h57ff3fff_00150184_2800018c_2600018c,
       128'h28ff62cc_29bfb2cc_02bf418c_0040818c,
       128'h001031ac_2800018c_270001cf_28ff62ce,
       128'h02c0058f_2600018c_28ff62cc_0040818d,
       128'h0040858c_0010358c_0040898c_001501ac,
       128'h28bfb2cd_50004400_29bfb2c0_29ff62c4,
       128'h02c0c076_29c08076_29c0a061_02ff4063,
       128'h4c000020_02c08063_28c06076_00150184,
       128'h0067818c_0340058c_0015000c_50000800,
       128'h0280040c_60000d8d_0280e40c_00005d8d,
       128'h2a3fbecc_64001d8d_0280bc0c_00005d8d,
       128'h2a3fbecc_293fbecc_0015008c_02c08076,
       128'h29c06076_02ff8063_4c000020_02c0c063,
       128'h28c0a076_00150184_0040818c_0011b1ac,
       128'h28ff62cc_28ffa2cd_47ffdd9f_29ff42cd,
       128'h02fffd8d_28ff42cc_40001580_2800018c,
       128'h28ffa2cc_29ffa2cc_02c0058c_28ffa2cc,
       128'h50001000_29ffa2cc_28ff62cc_29ff42c5,
       128'h29ff62c4_02c0c076_29c0a076_02ff4063,
       128'h4c000020_02c0c063_28c08076_28c0a061,
       128'h03400000_4c000181_001501a4_001501c5,
       128'h283fbecd_28c021ae_28ff82cd_2600018c,
       128'h28ff82cc_40002580_0067818c_2a3fbecc,
       128'h293fbecc_29ff42c7_29ff62c6_29ff82c5,
       128'h0015008c_02c0c076_29c08076_29c0a061,
       128'h02ff4063_4c000020_02c0c063_28c08076,
       128'h28c0a061_03400000_57fecbff_00150184,
       128'h283fbecc_40001180_0067818c_2a3fbecc,
       128'h293fbecc_29ff42c7_29ff62c6_29ff82c5,
       128'h0015008c_02c0c076_29c08076_29c0a061,
       128'h02ff4063_4c000020_02c0c063_28c0a076,
       128'h03400000_293fbecc_29ff42c7_29ff62c6,
       128'h29ff82c5_0015008c_02c0c076_29c0a076,
       128'h02ff4063_4c000020_02c0c063_28c0a076,
       128'h03400000_2900018d_2a3fbecd_0010b1ac,
       128'h28ff62cc_28ff82cd_6c0019ac_28ff42cc,
       128'h28ff62cd_293fbecc_29ff42c7_29ff62c6,
       128'h29ff82c5_0015008c_02c0c076_29c0a076,
       128'h02ff4063_4c000020_02c08063_28c04076,
       128'h28c06061_00150184_0015000c_57ff9fff,
       128'h00150184_00005d8c_28bfb2cc_29bfb2cc,
       128'h0015008c_02c08076_29c04076_29c06061,
       128'h02ff8063_4c000020_02c08063_28c04076,
       128'h28c06061_03400000_5428b000_00150184,
       128'h02bffc05_0040818c_283fbecc_293fbecc,
       128'h0015008c_02c08076_29c04076_29c06061,
       128'h02ff8063_4c000020_02c08063_28c04076,
       128'h28c06061_00150184_0015000c_5428f400,
       128'h02802804_02bffc05_47ffd99f_2800018c,
       128'h28ffa2cc_29ffa2cc_02c0058c_28ffa2cc,
       128'h54291800_00150184_02bffc05_2800018c,
       128'h28ffa2cc_50002400_29ffa2c4_02c08076,
       128'h29c04076_29c06061_02ff8063_4c000020,
       128'h02c0c063_28c0a076_00150184_24ffeecc,
       128'h63ffc9ac_0040818c_004081ad_28bf62cc,
       128'h28bfa2cd_29bfa2cc_001031ac_28bf52cc,
       128'h28bfa2cd_29bfb2cc_001031ac_28bfb2cd,
       128'h0040818c_0040858c_28bfa2cc_50002c00,
       128'h29bfa2c0_29bfb2cc_28bf72cc_29bf52cc,
       128'h001501ac_29bf62cc_001501cc_29bf72cc,
       128'h001500cd_001500ae_0015008c_02c0c076,
       128'h29c0a076_02ff4063_4c000020_02c14063,
       128'h28c10076_28c12061_00150184_0015000c,
       128'h5400a800_180157c4_5400b000_18015784,
       128'h48000c00_0c218400_0114a801_2bbec2c0,
       128'h54275400_18015784_28fee2c5_54276000,
       128'h18015764_28ff02c5_54276c00_18015744,
       128'h28ff22c5_54277800_18015724_28ff42c5,
       128'h54278400_18015704_28ff62c5_54279000,
       128'h180156e4_28ff82c5_29fec2c0_54011400,
       128'h18015664_2bfee2c0_01050020_2bbf02c0,
       128'h2bbf22c1_2bff02c0_01010020_2b800180,
       128'h18015cec_01050021_2b800180_18015e0c,
       128'h2bbfa2c1_2bff22c0_01010020_2b800180,
       128'h18015dec_01050021_2b800180_18015ecc,
       128'h2bbfa2c1_2bff42c0_01010020_2b800180,
       128'h18015eec_01050021_2b800180_18015f8c,
       128'h2bbfa2c1_2bff62c0_01010020_2b800180,
       128'h18015fec_01010001_2bbfa2c0_2bff82c0,
       128'h01010020_2b800180_180160ac_2bbfa2c1,
       128'h2bffa2c0_2b800180_180160ec_5401c400,
       128'h18015ae4_5401cc00_18015aa4_02c14076,
       128'h29c10076_29c12061_02fec063_54000000,
       128'h4c0000a0_38728000_38720000_29c000a4,
       128'h14a80004_180bf545_4c000181_0300018c,
       128'h1600000c_0385d18c_1438000c_01010421,
       128'h010304a5_011d2821_011d2061_011a8803,
       128'h38104188_38104188_38103d88_38103d88,
       128'h0380180f_38103987_38103987_0380140e,
       128'h0001b1a0_00013580_02c0198d_38103586,
       128'h38103585_03801c10_0380100d_0300018c,
       128'h1600000c_0380018c_1438008c_03840c08,
       128'h03844007_03840406_03840005_0400002c,
       128'h0380400c_0400082b_0380040b_0406042b,
       128'h0320016b_03803c0b_0406002b_0380440b,
       128'h28bfc2f8_030002f7_16000017_038002f7,
       128'h14380097_0015001f_0015001e_0015001d,
       128'h0015001c_0015001b_0015001a_00150019,
       128'h00150018_00150017_00150016_00150015,
       128'h00150014_00150013_00150012_00150011,
       128'h00150010_0015000f_0015000e_0015000d,
       128'h0015000c_0015000b_0015000a_00150009,
       128'h00150008_00150007_00150006_00150005,
       128'h00150004_03000063_16000003_03800063,
       128'h143800e3_00150002_00150001_4c000180,
       128'h0300018c_1600000c_0380518c_1438000c
};

/// read 
logic ram_cs;
// assign ram_cs = addr_i >= 64'h0000_0000 && addr_i < 64'h1FF0_0000;
assign ram_cs = addr_i[23:0] >= 24'h000000 && addr_i[23:0] < 24'hFFFFFF;
logic [AXI_ADDR_WIDTH-1:0] ram_raddr_q;
logic [AXI_DATA_WIDTH-1:0] ram_rdata_o;
always_ff @(posedge clk) begin
    if (ram_cs && req_i && ~ we_i) begin
        ram_raddr_q <= addr_i;
    end
end


logic [AXI_ADDR_WIDTH-1:0] ram_raddr; 

assign ram_raddr = ram_raddr_q[$clog2(RamSize)+3:4];
assign ram_rdata_o = reset ? '0 : ram_mem[ram_raddr];


/// write
logic [AXI_DATA_WIDTH-1:0] ram_rdata_i;

always_comb begin
    ram_rdata_i = ram_mem[addr_i[$clog2(RamSize)+3:4]];
    for (int i = 0; i < $bits(be_i); i++) begin
        if (be_i[i]) begin
            ram_rdata_i[i*8+:8] = data_i[i*8+:8];
        end
    end
end

always @(posedge clk) begin 
    if (ram_cs && req_i && we_i) begin
        ram_mem[addr_i[$clog2(RamSize)+3:4]] <= ram_rdata_i;
    end
end


/// --------------------------- UART --------------------------- ///

localparam int UARTSize = 1000;
logic [UARTSize-1:0][127:0] uart_map_mem = {
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000,
       128'h00000000_00000000_00000000_00000000
};

/// read 
logic UART_cs;
assign UART_cs = addr_i >= 64'h1FF1_0000 && addr_i < 64'h1FF1_FFFF;
logic [AXI_ADDR_WIDTH-1:0] UART_raddr_q;
logic [AXI_DATA_WIDTH-1:0] UART_rdata_o;
always_ff @(posedge clk) begin
    if (UART_cs && req_i && ~ we_i) begin
        UART_raddr_q <= addr_i;
    end
end
assign UART_rdata_o = (UART_raddr_q[AXI_ADDR_WIDTH-1:4] == 36'h1FF1_001) ? 128'h20_00000000 :
                      uart_map_mem[UART_raddr_q[$clog2(UARTSize)+3:4]];


/// write registers
logic [AXI_DATA_WIDTH-1:0] uart_rdata_i;

always_comb begin
    uart_rdata_i = uart_map_mem[addr_i[$clog2(RamSize)+3:4]];
    for (int i = 0; i < $bits(be_i); i++) begin
        if (be_i[i]) begin
            uart_rdata_i[i*8+:8] = data_i[i*8+:8];
        end
    end
end

always @(posedge clk) begin 
    if (UART_cs && req_i && we_i) begin
        uart_map_mem[addr_i[$clog2(RamSize)+3:4]] <= uart_rdata_i;
    end
end

/// write, print
always @(posedge clk) begin
     if (UART_cs && req_i && we_i) 
     begin
        if(be_i[15:0] == 16'h01) /// write 8-bit
           begin
              $write("%c", data_i[7:0]);
           end
        else if(be_i[15:0] == 16'hf) /// write 32-bit
           begin
              $write("%c", data_i[7:0]);
           end
        else if(be_i[15:0] == 16'hff) /// write 64-bit
           begin
              $write("%c", data_i[7:0]);
           end   
        else if(be_i[15:0] == 16'hf0)
           begin
              $write("%c", data_i[39:32]);
           end
        else if(be_i[15:0] == 16'hf00)
           begin
              $write("%c", data_i[71:64]);
           end
        else if(be_i[15:0] == 16'hf000)
           begin
              $write("%c", data_i[103:96]);
           end
    end
end

/// Read Data Output
always @(*) begin 
    if (ram_cs) begin
        data_o = ram_rdata_o;
    end
    else if (UART_cs) begin
        data_o = UART_rdata_o;
    end
    else begin
        data_o = '0;
    end
end

endmodule
